
module bch_encoder_p8 ( message, sel, code_o, clk, start, reset );
  input [7:0] message;
  output [7:0] code_o;
  input sel, clk, start, reset;
  wire   r0, r1, r2, r3, r4, r5, r6, r7, v8, v9, v10, v11, v12, v13, v14, v15,
         v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
         v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43,
         v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57,
         v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71,
         v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85,
         v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99,
         v100, v101, v102, v103, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571;
  wire   [7:0] message_r;
  wire   [7:0] parity;

  OAI222XL U2 ( .A0(n550), .A1(n3), .B0(n545), .B1(n5), .C0(n529), .C1(n7), 
        .Y(n391) );
  OAI222XL U3 ( .A0(n8), .A1(n9), .B0(v100), .B1(n10), .C0(n525), .C1(n11), 
        .Y(n392) );
  AOI22X1 U4 ( .A0(n521), .A1(n13), .B0(n516), .B1(n15), .Y(n10) );
  AOI221X1 U5 ( .A0(n14), .A1(n13), .B0(n12), .B1(n15), .C0(n538), .Y(n8) );
  OAI22X1 U6 ( .A0(n524), .A1(n9), .B0(n13), .B1(n549), .Y(n393) );
  INVX1 U7 ( .A(n15), .Y(n13) );
  INVX1 U8 ( .A(v100), .Y(n9) );
  OAI21XL U9 ( .A0(n6), .A1(n17), .B0(n18), .Y(n394) );
  AOI32X1 U10 ( .A0(n19), .A1(n20), .A2(n557), .B0(v102), .B1(n22), .Y(n18) );
  OAI22X1 U11 ( .A0(n524), .A1(n20), .B0(n23), .B1(n549), .Y(n395) );
  INVX1 U12 ( .A(v102), .Y(n20) );
  OAI222XL U13 ( .A0(n24), .A1(n25), .B0(v103), .B1(n26), .C0(n525), .C1(n27), 
        .Y(n396) );
  INVX1 U14 ( .A(v103), .Y(n25) );
  INVX1 U15 ( .A(n28), .Y(n397) );
  AOI222X1 U16 ( .A0(n29), .A1(n516), .B0(n30), .B1(n521), .C0(n536), .C1(v103), .Y(n28) );
  OAI21XL U17 ( .A0(n6), .A1(n32), .B0(n33), .Y(n398) );
  AOI32X1 U18 ( .A0(n34), .A1(n35), .A2(n556), .B0(v56), .B1(n36), .Y(n33) );
  OAI222XL U19 ( .A0(n37), .A1(n38), .B0(v64), .B1(n39), .C0(n525), .C1(n35), 
        .Y(n399) );
  INVX1 U20 ( .A(v56), .Y(n35) );
  AOI22X1 U21 ( .A0(n40), .A1(n12), .B0(n516), .B1(n41), .Y(n39) );
  AOI221X1 U22 ( .A0(n40), .A1(n14), .B0(n12), .B1(n41), .C0(n537), .Y(n37) );
  OAI21XL U23 ( .A0(n6), .A1(n38), .B0(n42), .Y(n400) );
  AOI32X1 U24 ( .A0(n43), .A1(n44), .A2(n556), .B0(v72), .B1(n45), .Y(n42) );
  OAI21XL U25 ( .A0(n551), .A1(n43), .B0(n541), .Y(n45) );
  INVX1 U26 ( .A(v64), .Y(n38) );
  OAI222XL U27 ( .A0(n46), .A1(n47), .B0(v80), .B1(n48), .C0(n525), .C1(n44), 
        .Y(n401) );
  INVX1 U28 ( .A(v72), .Y(n44) );
  AOI22X1 U29 ( .A0(n49), .A1(n521), .B0(n516), .B1(n50), .Y(n48) );
  AOI221X1 U30 ( .A0(n49), .A1(n14), .B0(n12), .B1(n50), .C0(n537), .Y(n46) );
  OAI222XL U31 ( .A0(n542), .A1(n51), .B0(n52), .B1(n553), .C0(n525), .C1(n47), 
        .Y(n402) );
  INVX1 U32 ( .A(v80), .Y(n47) );
  XNOR2X1 U33 ( .A(n53), .B(n54), .Y(n52) );
  XNOR2X1 U34 ( .A(v88), .B(n55), .Y(n53) );
  OAI222XL U35 ( .A0(n542), .A1(n56), .B0(n57), .B1(n552), .C0(n525), .C1(n58), 
        .Y(n403) );
  INVX1 U36 ( .A(v35), .Y(n58) );
  XOR2X1 U37 ( .A(n59), .B(n60), .Y(n57) );
  XNOR2X1 U38 ( .A(v43), .B(n34), .Y(n59) );
  OAI222XL U39 ( .A0(v51), .A1(n61), .B0(n62), .B1(n63), .C0(n525), .C1(n56), 
        .Y(n404) );
  INVX1 U40 ( .A(v43), .Y(n56) );
  AOI221X1 U41 ( .A0(n64), .A1(n65), .B0(n66), .B1(n67), .C0(n537), .Y(n62) );
  OAI21XL U42 ( .A0(n534), .A1(n63), .B0(n68), .Y(n405) );
  AOI32X1 U43 ( .A0(n69), .A1(n70), .A2(n556), .B0(v59), .B1(n71), .Y(n68) );
  INVX1 U44 ( .A(v51), .Y(n63) );
  OAI222XL U45 ( .A0(n72), .A1(n73), .B0(v67), .B1(n74), .C0(n525), .C1(n70), 
        .Y(n406) );
  INVX1 U46 ( .A(v59), .Y(n70) );
  AOI22X1 U47 ( .A0(n75), .A1(n76), .B0(n77), .B1(n78), .Y(n74) );
  AOI221X1 U48 ( .A0(n77), .A1(n76), .B0(n75), .B1(n78), .C0(n537), .Y(n72) );
  OAI222XL U49 ( .A0(n79), .A1(n80), .B0(v75), .B1(n81), .C0(n525), .C1(n73), 
        .Y(n407) );
  INVX1 U50 ( .A(v67), .Y(n73) );
  OAI222XL U51 ( .A0(n82), .A1(n83), .B0(v83), .B1(n84), .C0(n526), .C1(n80), 
        .Y(n408) );
  INVX1 U52 ( .A(v75), .Y(n80) );
  AOI22X1 U53 ( .A0(n85), .A1(n66), .B0(n64), .B1(n86), .Y(n84) );
  AOI221X1 U54 ( .A0(n85), .A1(n64), .B0(n66), .B1(n86), .C0(n537), .Y(n82) );
  OAI21XL U55 ( .A0(n534), .A1(n83), .B0(n87), .Y(n409) );
  AOI32X1 U56 ( .A0(n88), .A1(n89), .A2(n523), .B0(v91), .B1(n90), .Y(n87) );
  INVX1 U57 ( .A(v83), .Y(n83) );
  OAI222XL U58 ( .A0(n91), .A1(n92), .B0(v99), .B1(n93), .C0(n526), .C1(n89), 
        .Y(n410) );
  INVX1 U59 ( .A(v91), .Y(n89) );
  AOI22X1 U60 ( .A0(n518), .A1(n95), .B0(n522), .B1(n19), .Y(n93) );
  AOI221X1 U61 ( .A0(n94), .A1(n19), .B0(n96), .B1(n95), .C0(n537), .Y(n91) );
  INVX1 U62 ( .A(n19), .Y(n95) );
  OAI21XL U63 ( .A0(n533), .A1(n92), .B0(n97), .Y(n411) );
  INVX1 U64 ( .A(v99), .Y(n92) );
  OAI222XL U65 ( .A0(n550), .A1(n98), .B0(n544), .B1(n99), .C0(n526), .C1(n100), .Y(n412) );
  OAI222XL U66 ( .A0(n542), .A1(n101), .B0(n102), .B1(n553), .C0(n526), .C1(
        n99), .Y(n413) );
  XOR2X1 U67 ( .A(n103), .B(n104), .Y(n102) );
  XNOR2X1 U68 ( .A(v11), .B(n105), .Y(n103) );
  OAI21XL U69 ( .A0(n534), .A1(n101), .B0(n106), .Y(n414) );
  AOI32X1 U70 ( .A0(n19), .A1(n107), .A2(n523), .B0(v19), .B1(n22), .Y(n106)
         );
  OAI21XL U71 ( .A0(n551), .A1(n19), .B0(n542), .Y(n22) );
  XNOR2X1 U72 ( .A(n108), .B(n65), .Y(n19) );
  INVX1 U73 ( .A(v11), .Y(n101) );
  OAI222XL U74 ( .A0(n109), .A1(n110), .B0(v27), .B1(n111), .C0(n526), .C1(
        n107), .Y(n415) );
  INVX1 U75 ( .A(v19), .Y(n107) );
  AOI22X1 U76 ( .A0(n512), .A1(n113), .B0(n513), .B1(n115), .Y(n111) );
  AOI221X1 U77 ( .A0(n112), .A1(n115), .B0(n114), .B1(n113), .C0(n537), .Y(
        n109) );
  OAI22X1 U78 ( .A0(n54), .A1(n116), .B0(n117), .B1(n118), .Y(n113) );
  OAI22X1 U79 ( .A0(n117), .A1(n116), .B0(n54), .B1(n118), .Y(n115) );
  INVX1 U80 ( .A(n117), .Y(n54) );
  OAI221XL U81 ( .A0(v35), .A1(n119), .B0(n532), .B1(n110), .C0(n120), .Y(n416) );
  OAI21XL U82 ( .A0(n121), .A1(n540), .B0(v35), .Y(n120) );
  INVX1 U83 ( .A(v27), .Y(n110) );
  OAI222XL U84 ( .A0(n543), .A1(n122), .B0(n123), .B1(n552), .C0(n526), .C1(
        n51), .Y(n417) );
  INVX1 U85 ( .A(v88), .Y(n51) );
  XOR2X1 U86 ( .A(n124), .B(n125), .Y(n123) );
  XNOR2X1 U87 ( .A(v96), .B(n67), .Y(n124) );
  OAI222XL U88 ( .A0(n543), .A1(n126), .B0(n127), .B1(n553), .C0(n526), .C1(
        n128), .Y(n418) );
  XNOR2X1 U89 ( .A(n104), .B(n129), .Y(n127) );
  XNOR2X1 U90 ( .A(n126), .B(n55), .Y(n129) );
  OAI21XL U91 ( .A0(n533), .A1(n126), .B0(n61), .Y(n419) );
  AOI22X1 U92 ( .A0(n67), .A1(n64), .B0(n65), .B1(n66), .Y(n61) );
  INVX1 U93 ( .A(v101), .Y(n126) );
  OAI22X1 U94 ( .A0(n525), .A1(n122), .B0(n130), .B1(n549), .Y(n420) );
  INVX1 U95 ( .A(v96), .Y(n122) );
  OAI222XL U96 ( .A0(n550), .A1(n131), .B0(n545), .B1(n132), .C0(n526), .C1(
        n133), .Y(n421) );
  OAI222XL U97 ( .A0(n134), .A1(n135), .B0(v8), .B1(n136), .C0(n526), .C1(n132), .Y(n422) );
  AOI22X1 U98 ( .A0(n522), .A1(n513), .B0(n518), .B1(n112), .Y(n136) );
  AOI221X1 U99 ( .A0(n94), .A1(n114), .B0(n96), .B1(n112), .C0(n537), .Y(n134)
         );
  OAI222XL U100 ( .A0(n544), .A1(n137), .B0(n138), .B1(n553), .C0(n526), .C1(
        n135), .Y(n423) );
  INVX1 U101 ( .A(v8), .Y(n135) );
  XNOR2X1 U102 ( .A(n139), .B(n140), .Y(n138) );
  XNOR2X1 U103 ( .A(v16), .B(n141), .Y(n139) );
  OAI222XL U104 ( .A0(n142), .A1(n143), .B0(v24), .B1(n144), .C0(n527), .C1(
        n137), .Y(n424) );
  INVX1 U105 ( .A(v16), .Y(n137) );
  AOI22X1 U106 ( .A0(n522), .A1(n41), .B0(n518), .B1(n40), .Y(n144) );
  AOI221X1 U107 ( .A0(n518), .A1(n41), .B0(n96), .B1(n40), .C0(n537), .Y(n142)
         );
  INVX1 U108 ( .A(n41), .Y(n40) );
  XNOR2X1 U109 ( .A(n145), .B(n112), .Y(n41) );
  OAI222XL U110 ( .A0(n543), .A1(n146), .B0(n147), .B1(n553), .C0(n527), .C1(
        n143), .Y(n425) );
  INVX1 U111 ( .A(v24), .Y(n143) );
  XNOR2X1 U112 ( .A(n148), .B(n149), .Y(n147) );
  XNOR2X1 U113 ( .A(v32), .B(n150), .Y(n148) );
  OAI222XL U114 ( .A0(n544), .A1(n151), .B0(n152), .B1(n553), .C0(n527), .C1(
        n146), .Y(n426) );
  INVX1 U115 ( .A(v32), .Y(n146) );
  XNOR2X1 U116 ( .A(n153), .B(n140), .Y(n152) );
  XNOR2X1 U117 ( .A(v40), .B(n78), .Y(n153) );
  OAI21XL U118 ( .A0(n534), .A1(n151), .B0(n154), .Y(n427) );
  AOI32X1 U119 ( .A0(n515), .A1(n32), .A2(n523), .B0(v48), .B1(n155), .Y(n154)
         );
  OAI21XL U120 ( .A0(n552), .A1(n86), .B0(n4), .Y(n155) );
  INVX1 U121 ( .A(v48), .Y(n32) );
  INVX1 U122 ( .A(v40), .Y(n151) );
  OAI222XL U123 ( .A0(n551), .A1(n156), .B0(n545), .B1(n157), .C0(n527), .C1(
        n158), .Y(n428) );
  OAI222XL U124 ( .A0(n544), .A1(n159), .B0(n160), .B1(n553), .C0(n527), .C1(
        n157), .Y(n429) );
  XOR2X1 U125 ( .A(n161), .B(n162), .Y(n160) );
  XNOR2X1 U126 ( .A(v10), .B(n55), .Y(n161) );
  OAI222XL U127 ( .A0(n163), .A1(n164), .B0(v18), .B1(n165), .C0(n527), .C1(
        n159), .Y(n430) );
  INVX1 U128 ( .A(v10), .Y(n159) );
  AOI22X1 U129 ( .A0(n166), .A1(n521), .B0(n516), .B1(n167), .Y(n165) );
  AOI221X1 U130 ( .A0(n166), .A1(n14), .B0(n12), .B1(n167), .C0(n538), .Y(n163) );
  INVX1 U131 ( .A(n167), .Y(n166) );
  OAI222XL U132 ( .A0(n168), .A1(n169), .B0(v26), .B1(n170), .C0(n527), .C1(
        n164), .Y(n431) );
  INVX1 U133 ( .A(v18), .Y(n164) );
  AOI22X1 U134 ( .A0(n522), .A1(n67), .B0(n518), .B1(n65), .Y(n170) );
  AOI221X1 U135 ( .A0(n94), .A1(n67), .B0(n96), .B1(n65), .C0(n538), .Y(n168)
         );
  OAI21XL U136 ( .A0(n534), .A1(n169), .B0(n171), .Y(n432) );
  AOI32X1 U137 ( .A0(n117), .A1(n172), .A2(n523), .B0(v34), .B1(n173), .Y(n171) );
  OAI21XL U138 ( .A0(n552), .A1(n117), .B0(n4), .Y(n173) );
  XOR2X1 U139 ( .A(n174), .B(n175), .Y(n117) );
  INVX1 U140 ( .A(v26), .Y(n169) );
  OAI21XL U141 ( .A0(n533), .A1(n172), .B0(n176), .Y(n433) );
  AOI32X1 U142 ( .A0(n177), .A1(n178), .A2(n523), .B0(v42), .B1(n179), .Y(n176) );
  INVX1 U143 ( .A(v34), .Y(n172) );
  OAI21XL U144 ( .A0(n533), .A1(n178), .B0(n180), .Y(n434) );
  AOI32X1 U145 ( .A0(n15), .A1(n181), .A2(n523), .B0(v50), .B1(n182), .Y(n180)
         );
  OAI21XL U146 ( .A0(n552), .A1(n15), .B0(n545), .Y(n182) );
  INVX1 U147 ( .A(v42), .Y(n178) );
  OAI222XL U148 ( .A0(n183), .A1(n184), .B0(v58), .B1(n185), .C0(n527), .C1(
        n181), .Y(n435) );
  INVX1 U149 ( .A(v50), .Y(n181) );
  OAI222XL U150 ( .A0(n186), .A1(n187), .B0(v66), .B1(n188), .C0(n527), .C1(
        n184), .Y(n436) );
  INVX1 U151 ( .A(v58), .Y(n184) );
  AOI22X1 U152 ( .A0(n522), .A1(n515), .B0(n518), .B1(n85), .Y(n188) );
  AOI221X1 U153 ( .A0(n94), .A1(n86), .B0(n96), .B1(n85), .C0(n538), .Y(n186)
         );
  OAI222XL U154 ( .A0(n189), .A1(n190), .B0(v74), .B1(n191), .C0(n527), .C1(
        n187), .Y(n437) );
  INVX1 U155 ( .A(v66), .Y(n187) );
  OAI222XL U156 ( .A0(n544), .A1(n192), .B0(n193), .B1(n553), .C0(n528), .C1(
        n190), .Y(n438) );
  INVX1 U157 ( .A(v74), .Y(n190) );
  XNOR2X1 U158 ( .A(n194), .B(n195), .Y(n193) );
  XNOR2X1 U159 ( .A(v82), .B(n114), .Y(n194) );
  OAI21XL U160 ( .A0(n533), .A1(n192), .B0(n196), .Y(n439) );
  AOI32X1 U161 ( .A0(n34), .A1(n197), .A2(n523), .B0(v90), .B1(n36), .Y(n196)
         );
  OAI21XL U162 ( .A0(n552), .A1(n34), .B0(n545), .Y(n36) );
  INVX1 U163 ( .A(v82), .Y(n192) );
  OAI21XL U164 ( .A0(n534), .A1(n197), .B0(n198), .Y(n440) );
  AOI32X1 U165 ( .A0(n177), .A1(n199), .A2(n555), .B0(v98), .B1(n179), .Y(n198) );
  OAI21XL U166 ( .A0(n552), .A1(n177), .B0(n545), .Y(n179) );
  INVX1 U167 ( .A(v98), .Y(n199) );
  XNOR2X1 U168 ( .A(n200), .B(n167), .Y(n177) );
  XNOR2X1 U169 ( .A(n55), .B(n130), .Y(n167) );
  INVX1 U170 ( .A(v90), .Y(n197) );
  INVX1 U171 ( .A(n201), .Y(n441) );
  AOI222X1 U172 ( .A0(n105), .A1(n202), .B0(n203), .B1(n204), .C0(n536), .C1(
        v98), .Y(n201) );
  OAI222XL U173 ( .A0(n550), .A1(n205), .B0(n545), .B1(n206), .C0(n528), .C1(
        n207), .Y(n442) );
  OAI222XL U174 ( .A0(n544), .A1(n208), .B0(n209), .B1(n553), .C0(n528), .C1(
        n206), .Y(n443) );
  XNOR2X1 U175 ( .A(n125), .B(n210), .Y(n209) );
  XNOR2X1 U176 ( .A(n208), .B(n55), .Y(n210) );
  OAI21XL U177 ( .A0(n533), .A1(n208), .B0(n211), .Y(n444) );
  AOI32X1 U178 ( .A0(n108), .A1(n212), .A2(n555), .B0(v23), .B1(n213), .Y(n211) );
  OAI21XL U179 ( .A0(n552), .A1(n108), .B0(n4), .Y(n213) );
  INVX1 U180 ( .A(v15), .Y(n208) );
  OAI222XL U181 ( .A0(n214), .A1(n215), .B0(v31), .B1(n216), .C0(n528), .C1(
        n212), .Y(n445) );
  INVX1 U182 ( .A(v23), .Y(n212) );
  OAI222XL U183 ( .A0(n544), .A1(n217), .B0(n218), .B1(n554), .C0(n528), .C1(
        n215), .Y(n446) );
  INVX1 U184 ( .A(v31), .Y(n215) );
  XOR2X1 U185 ( .A(n219), .B(n220), .Y(n218) );
  XNOR2X1 U186 ( .A(v39), .B(n86), .Y(n219) );
  OAI222XL U187 ( .A0(n221), .A1(n222), .B0(v47), .B1(n223), .C0(n528), .C1(
        n217), .Y(n447) );
  INVX1 U188 ( .A(v39), .Y(n217) );
  AOI22X1 U189 ( .A0(n512), .A1(n521), .B0(n14), .B1(n114), .Y(n223) );
  AOI221X1 U190 ( .A0(n112), .A1(n14), .B0(n12), .B1(n114), .C0(n538), .Y(n221) );
  OAI21XL U191 ( .A0(n534), .A1(n222), .B0(n224), .Y(n448) );
  AOI32X1 U192 ( .A0(n78), .A1(n225), .A2(n557), .B0(v55), .B1(n226), .Y(n224)
         );
  OAI21XL U193 ( .A0(n552), .A1(n78), .B0(n4), .Y(n226) );
  INVX1 U194 ( .A(v47), .Y(n222) );
  OAI21XL U195 ( .A0(n534), .A1(n225), .B0(n227), .Y(n449) );
  AOI32X1 U196 ( .A0(n228), .A1(n229), .A2(n523), .B0(v63), .B1(n230), .Y(n227) );
  INVX1 U197 ( .A(v55), .Y(n225) );
  OAI222XL U198 ( .A0(n231), .A1(n232), .B0(v71), .B1(n233), .C0(n528), .C1(
        n229), .Y(n450) );
  INVX1 U199 ( .A(v63), .Y(n229) );
  AOI22X1 U200 ( .A0(n66), .A1(n234), .B0(n520), .B1(n174), .Y(n233) );
  AOI221X1 U201 ( .A0(n64), .A1(n234), .B0(n66), .B1(n174), .C0(n538), .Y(n231) );
  OAI222XL U202 ( .A0(n235), .A1(n236), .B0(v79), .B1(n237), .C0(n528), .C1(
        n232), .Y(n451) );
  INVX1 U203 ( .A(v71), .Y(n232) );
  OAI222XL U204 ( .A0(n235), .A1(n238), .B0(v87), .B1(n237), .C0(n528), .C1(
        n236), .Y(n452) );
  INVX1 U205 ( .A(v79), .Y(n236) );
  AOI22X1 U206 ( .A0(n239), .A1(n64), .B0(n66), .B1(n23), .Y(n237) );
  AOI221X1 U207 ( .A0(n239), .A1(n517), .B0(n64), .B1(n23), .C0(n538), .Y(n235) );
  INVX1 U208 ( .A(n239), .Y(n23) );
  OAI222XL U209 ( .A0(n544), .A1(n27), .B0(n240), .B1(n554), .C0(n528), .C1(
        n238), .Y(n453) );
  INVX1 U210 ( .A(v87), .Y(n238) );
  XNOR2X1 U211 ( .A(n241), .B(n242), .Y(n240) );
  XNOR2X1 U212 ( .A(v95), .B(n15), .Y(n241) );
  INVX1 U213 ( .A(v95), .Y(n27) );
  OAI222XL U214 ( .A0(n550), .A1(n243), .B0(n545), .B1(n244), .C0(n529), .C1(
        n245), .Y(n454) );
  OAI222XL U215 ( .A0(n246), .A1(n247), .B0(v14), .B1(n248), .C0(n529), .C1(
        n244), .Y(n455) );
  AOI22X1 U216 ( .A0(n242), .A1(n75), .B0(n77), .B1(n249), .Y(n248) );
  AOI221X1 U217 ( .A0(n242), .A1(n77), .B0(n75), .B1(n249), .C0(n538), .Y(n246) );
  OAI21XL U218 ( .A0(n533), .A1(n247), .B0(n250), .Y(n456) );
  AOI32X1 U219 ( .A0(n55), .A1(n251), .A2(n555), .B0(v22), .B1(n252), .Y(n250)
         );
  OAI21XL U220 ( .A0(n551), .A1(n55), .B0(n541), .Y(n252) );
  INVX1 U221 ( .A(v14), .Y(n247) );
  OAI222XL U222 ( .A0(n253), .A1(n254), .B0(v30), .B1(n255), .C0(n529), .C1(
        n251), .Y(n457) );
  INVX1 U223 ( .A(v22), .Y(n251) );
  OAI222XL U224 ( .A0(n544), .A1(n256), .B0(n257), .B1(n554), .C0(n529), .C1(
        n254), .Y(n458) );
  INVX1 U225 ( .A(v30), .Y(n254) );
  XNOR2X1 U226 ( .A(n258), .B(n85), .Y(n257) );
  XNOR2X1 U227 ( .A(v38), .B(n162), .Y(n258) );
  OAI21XL U228 ( .A0(n533), .A1(n256), .B0(n259), .Y(n459) );
  AOI32X1 U229 ( .A0(n228), .A1(n260), .A2(n555), .B0(v46), .B1(n230), .Y(n259) );
  OAI21XL U230 ( .A0(n551), .A1(n228), .B0(n542), .Y(n230) );
  INVX1 U231 ( .A(v38), .Y(n256) );
  OAI21XL U232 ( .A0(n533), .A1(n260), .B0(n261), .Y(n460) );
  AOI32X1 U233 ( .A0(n513), .A1(n262), .A2(n557), .B0(v54), .B1(n263), .Y(n261) );
  OAI21XL U234 ( .A0(n551), .A1(n513), .B0(n4), .Y(n263) );
  INVX1 U235 ( .A(v46), .Y(n260) );
  OAI222XL U236 ( .A0(n264), .A1(n265), .B0(v62), .B1(n266), .C0(n529), .C1(
        n262), .Y(n461) );
  INVX1 U237 ( .A(v54), .Y(n262) );
  AOI22X1 U238 ( .A0(n149), .A1(n66), .B0(n64), .B1(n228), .Y(n266) );
  AOI221X1 U239 ( .A0(n149), .A1(n64), .B0(n66), .B1(n228), .C0(n538), .Y(n264) );
  OAI222XL U240 ( .A0(n543), .A1(n267), .B0(n268), .B1(n554), .C0(n529), .C1(
        n265), .Y(n462) );
  INVX1 U241 ( .A(v62), .Y(n265) );
  XNOR2X1 U242 ( .A(n269), .B(n149), .Y(n268) );
  XNOR2X1 U243 ( .A(v70), .B(n34), .Y(n269) );
  OAI222XL U244 ( .A0(n270), .A1(n271), .B0(v78), .B1(n272), .C0(n530), .C1(
        n267), .Y(n463) );
  INVX1 U245 ( .A(v70), .Y(n267) );
  OAI222XL U246 ( .A0(n270), .A1(n273), .B0(v86), .B1(n272), .C0(n529), .C1(
        n271), .Y(n464) );
  INVX1 U247 ( .A(v78), .Y(n271) );
  AOI22X1 U248 ( .A0(n67), .A1(n77), .B0(n65), .B1(n75), .Y(n272) );
  AOI221X1 U249 ( .A0(n67), .A1(n75), .B0(n65), .B1(n77), .C0(n538), .Y(n270)
         );
  OAI222XL U250 ( .A0(n274), .A1(n17), .B0(v94), .B1(n275), .C0(n529), .C1(
        n273), .Y(n465) );
  INVX1 U251 ( .A(v86), .Y(n273) );
  AOI22X1 U252 ( .A0(n276), .A1(n75), .B0(n77), .B1(n277), .Y(n275) );
  INVX1 U253 ( .A(v94), .Y(n17) );
  AOI221X1 U254 ( .A0(n276), .A1(n77), .B0(n75), .B1(n277), .C0(n539), .Y(n274) );
  OAI222XL U255 ( .A0(n543), .A1(n278), .B0(n279), .B1(n554), .C0(n5), .C1(
        n533), .Y(n466) );
  XOR2X1 U256 ( .A(n280), .B(n220), .Y(n279) );
  XNOR2X1 U257 ( .A(v13), .B(n105), .Y(n280) );
  OAI221XL U258 ( .A0(v21), .A1(n118), .B0(n532), .B1(n278), .C0(n281), .Y(
        n467) );
  OAI21XL U259 ( .A0(n520), .A1(n540), .B0(v21), .Y(n281) );
  INVX1 U260 ( .A(v13), .Y(n278) );
  OAI2BB1X1 U261 ( .A0N(n535), .A1N(v21), .B0(n282), .Y(n468) );
  AOI32X1 U262 ( .A0(n69), .A1(n283), .A2(n557), .B0(v29), .B1(n71), .Y(n282)
         );
  OAI21XL U263 ( .A0(n551), .A1(n69), .B0(n542), .Y(n71) );
  XNOR2X1 U264 ( .A(n203), .B(n162), .Y(n69) );
  OAI222XL U265 ( .A0(n284), .A1(n285), .B0(v37), .B1(n286), .C0(n530), .C1(
        n283), .Y(n469) );
  INVX1 U266 ( .A(v29), .Y(n283) );
  AOI22X1 U267 ( .A0(n121), .A1(n86), .B0(n287), .B1(n85), .Y(n286) );
  AOI221X1 U268 ( .A0(n287), .A1(n86), .B0(n121), .B1(n85), .C0(n539), .Y(n284) );
  OAI222XL U269 ( .A0(n288), .A1(n289), .B0(v45), .B1(n290), .C0(n530), .C1(
        n285), .Y(n470) );
  INVX1 U270 ( .A(v37), .Y(n285) );
  AOI22X1 U271 ( .A0(n30), .A1(n291), .B0(n29), .B1(n292), .Y(n290) );
  AOI221X1 U272 ( .A0(n30), .A1(n292), .B0(n29), .B1(n291), .C0(n539), .Y(n288) );
  OAI22X1 U273 ( .A0(n293), .A1(n116), .B0(n43), .B1(n118), .Y(n291) );
  OAI22X1 U274 ( .A0(n43), .A1(n116), .B0(n293), .B1(n118), .Y(n292) );
  INVX1 U275 ( .A(n66), .Y(n118) );
  INVX1 U277 ( .A(n64), .Y(n116) );
  OAI221XL U279 ( .A0(v53), .A1(n296), .B0(n532), .B1(n289), .C0(n297), .Y(
        n471) );
  OAI21XL U280 ( .A0(n516), .A1(n540), .B0(v53), .Y(n297) );
  INVX1 U281 ( .A(v45), .Y(n289) );
  INVX1 U282 ( .A(n12), .Y(n296) );
  OAI222XL U283 ( .A0(n214), .A1(n298), .B0(v61), .B1(n216), .C0(n531), .C1(
        n299), .Y(n472) );
  INVX1 U284 ( .A(v53), .Y(n299) );
  AOI22X1 U285 ( .A0(n300), .A1(n202), .B0(n204), .B1(n140), .Y(n216) );
  AOI221X1 U286 ( .A0(n300), .A1(n204), .B0(n202), .B1(n140), .C0(n539), .Y(
        n214) );
  INVX1 U287 ( .A(n300), .Y(n140) );
  XNOR2X1 U288 ( .A(n43), .B(n301), .Y(n300) );
  OAI222XL U289 ( .A0(n543), .A1(n302), .B0(n303), .B1(n554), .C0(n530), .C1(
        n298), .Y(n473) );
  INVX1 U290 ( .A(v61), .Y(n298) );
  XNOR2X1 U291 ( .A(n304), .B(n130), .Y(n303) );
  XNOR2X1 U292 ( .A(v69), .B(n60), .Y(n304) );
  XNOR2X1 U293 ( .A(n293), .B(n108), .Y(n60) );
  INVX1 U294 ( .A(n43), .Y(n293) );
  OAI222XL U295 ( .A0(n253), .A1(n305), .B0(v77), .B1(n255), .C0(n531), .C1(
        n302), .Y(n474) );
  INVX1 U296 ( .A(v69), .Y(n302) );
  OAI222XL U297 ( .A0(n543), .A1(n306), .B0(n307), .B1(n554), .C0(n530), .C1(
        n305), .Y(n475) );
  INVX1 U298 ( .A(v77), .Y(n305) );
  XNOR2X1 U299 ( .A(n125), .B(n308), .Y(n307) );
  XNOR2X1 U300 ( .A(n306), .B(n145), .Y(n308) );
  XOR2X1 U301 ( .A(n108), .B(n309), .Y(n125) );
  OAI222XL U302 ( .A0(n310), .A1(n128), .B0(v93), .B1(n311), .C0(n530), .C1(
        n306), .Y(n476) );
  INVX1 U303 ( .A(v85), .Y(n306) );
  AOI22X1 U304 ( .A0(n522), .A1(n105), .B0(n518), .B1(n203), .Y(n311) );
  INVX1 U305 ( .A(v93), .Y(n128) );
  AOI221X1 U306 ( .A0(n94), .A1(n105), .B0(n96), .B1(n203), .C0(n539), .Y(n310) );
  INVX1 U307 ( .A(n105), .Y(n203) );
  XNOR2X1 U308 ( .A(n108), .B(n112), .Y(n105) );
  OAI222XL U309 ( .A0(n550), .A1(n312), .B0(n545), .B1(n313), .C0(n531), .C1(
        n314), .Y(n477) );
  OAI222XL U310 ( .A0(n543), .A1(n315), .B0(n316), .B1(n554), .C0(n530), .C1(
        n313), .Y(n478) );
  XNOR2X1 U311 ( .A(n317), .B(n242), .Y(n316) );
  XNOR2X1 U312 ( .A(v12), .B(n162), .Y(n317) );
  XNOR2X1 U313 ( .A(n318), .B(n175), .Y(n162) );
  OAI222XL U314 ( .A0(n24), .A1(n319), .B0(v20), .B1(n26), .C0(n531), .C1(n315), .Y(n479) );
  INVX1 U315 ( .A(v12), .Y(n315) );
  AOI22X1 U316 ( .A0(n34), .A1(n14), .B0(n12), .B1(n195), .Y(n26) );
  AOI221X1 U317 ( .A0(n34), .A1(n12), .B0(n14), .B1(n195), .C0(n539), .Y(n24)
         );
  INVX1 U318 ( .A(n34), .Y(n195) );
  XNOR2X1 U319 ( .A(n320), .B(n30), .Y(n34) );
  OAI222XL U320 ( .A0(n183), .A1(n321), .B0(v28), .B1(n185), .C0(n530), .C1(
        n319), .Y(n480) );
  INVX1 U321 ( .A(v20), .Y(n319) );
  AOI22X1 U322 ( .A0(n287), .A1(n242), .B0(n249), .B1(n121), .Y(n185) );
  AOI221X1 U323 ( .A0(n121), .A1(n514), .B0(n249), .B1(n287), .C0(n539), .Y(
        n183) );
  OAI222XL U324 ( .A0(n189), .A1(n322), .B0(v36), .B1(n191), .C0(n532), .C1(
        n321), .Y(n481) );
  INVX1 U325 ( .A(v28), .Y(n321) );
  AOI22X1 U326 ( .A0(n112), .A1(n287), .B0(n114), .B1(n121), .Y(n191) );
  AOI221X1 U327 ( .A0(n112), .A1(n121), .B0(n114), .B1(n287), .C0(n539), .Y(
        n189) );
  OAI222XL U328 ( .A0(n543), .A1(n323), .B0(n324), .B1(n554), .C0(n529), .C1(
        n322), .Y(n482) );
  INVX1 U329 ( .A(v36), .Y(n322) );
  XOR2X1 U330 ( .A(n325), .B(n326), .Y(n324) );
  XNOR2X1 U331 ( .A(n323), .B(n145), .Y(n326) );
  OAI222XL U332 ( .A0(n327), .A1(n328), .B0(v52), .B1(n329), .C0(n531), .C1(
        n323), .Y(n483) );
  INVX1 U333 ( .A(v44), .Y(n323) );
  AOI22X1 U334 ( .A0(n149), .A1(n204), .B0(n202), .B1(n228), .Y(n329) );
  AOI221X1 U335 ( .A0(n149), .A1(n202), .B0(n204), .B1(n228), .C0(n539), .Y(
        n327) );
  INVX1 U336 ( .A(n228), .Y(n149) );
  OAI222XL U337 ( .A0(n253), .A1(n330), .B0(v60), .B1(n255), .C0(n530), .C1(
        n328), .Y(n484) );
  INVX1 U338 ( .A(v52), .Y(n328) );
  NAND2X1 U339 ( .A(n557), .B(n331), .Y(n255) );
  AOI2BB1X1 U340 ( .A0N(n547), .A1N(n331), .B0(n540), .Y(n253) );
  XOR2X1 U341 ( .A(n332), .B(n15), .Y(n331) );
  XOR2X1 U342 ( .A(n309), .B(n175), .Y(n15) );
  OAI222XL U343 ( .A0(n333), .A1(n334), .B0(v68), .B1(n335), .C0(n532), .C1(
        n330), .Y(n485) );
  INVX1 U344 ( .A(v60), .Y(n330) );
  AOI22X1 U345 ( .A0(n75), .A1(n49), .B0(n77), .B1(n50), .Y(n335) );
  AOI221X1 U346 ( .A0(n77), .A1(n49), .B0(n75), .B1(n50), .C0(n540), .Y(n333)
         );
  INVX1 U348 ( .A(n309), .Y(n301) );
  INVX1 U349 ( .A(n50), .Y(n49) );
  OAI222XL U351 ( .A0(n336), .A1(n337), .B0(v76), .B1(n338), .C0(n532), .C1(
        n334), .Y(n486) );
  INVX1 U352 ( .A(v68), .Y(n334) );
  AOI22X1 U353 ( .A0(n522), .A1(n277), .B0(n276), .B1(n518), .Y(n338) );
  AOI221X1 U354 ( .A0(n94), .A1(n277), .B0(n276), .B1(n96), .C0(n540), .Y(n336) );
  INVX1 U355 ( .A(n277), .Y(n276) );
  XNOR2X1 U356 ( .A(n145), .B(n511), .Y(n277) );
  OAI222XL U357 ( .A0(n339), .A1(n340), .B0(v84), .B1(n341), .C0(n531), .C1(
        n337), .Y(n487) );
  INVX1 U358 ( .A(v76), .Y(n337) );
  AOI22X1 U359 ( .A0(n522), .A1(n249), .B0(n242), .B1(n518), .Y(n341) );
  AOI221X1 U360 ( .A0(n94), .A1(n249), .B0(n242), .B1(n96), .C0(n540), .Y(n339) );
  OAI222XL U361 ( .A0(n342), .A1(n11), .B0(v92), .B1(n343), .C0(n531), .C1(
        n340), .Y(n488) );
  INVX1 U362 ( .A(v84), .Y(n340) );
  AOI22X1 U363 ( .A0(n242), .A1(n204), .B0(n202), .B1(n249), .Y(n343) );
  INVX1 U364 ( .A(v92), .Y(n11) );
  AOI221X1 U365 ( .A0(n242), .A1(n202), .B0(n204), .B1(n249), .C0(n540), .Y(
        n342) );
  INVX1 U366 ( .A(n242), .Y(n249) );
  OAI222XL U368 ( .A0(n550), .A1(n345), .B0(n545), .B1(n346), .C0(n531), .C1(
        n347), .Y(n489) );
  OAI222XL U369 ( .A0(n542), .A1(n348), .B0(n349), .B1(n547), .C0(n531), .C1(
        n346), .Y(n490) );
  XNOR2X1 U370 ( .A(n350), .B(n130), .Y(n349) );
  XNOR2X1 U371 ( .A(v9), .B(n332), .Y(n350) );
  OAI222XL U372 ( .A0(n542), .A1(n351), .B0(n352), .B1(n554), .C0(n531), .C1(
        n348), .Y(n491) );
  INVX1 U373 ( .A(v9), .Y(n348) );
  XOR2X1 U374 ( .A(n353), .B(n220), .Y(n352) );
  XNOR2X1 U375 ( .A(n30), .B(n309), .Y(n220) );
  XNOR2X1 U376 ( .A(v17), .B(n228), .Y(n353) );
  OAI222XL U378 ( .A0(n542), .A1(n354), .B0(n355), .B1(n553), .C0(n530), .C1(
        n351), .Y(n492) );
  INVX1 U379 ( .A(v17), .Y(n351) );
  XNOR2X1 U380 ( .A(n104), .B(n356), .Y(n355) );
  XNOR2X1 U381 ( .A(n354), .B(n332), .Y(n356) );
  XOR2X1 U382 ( .A(n295), .B(n175), .Y(n104) );
  OAI21XL U383 ( .A0(n534), .A1(n354), .B0(n357), .Y(n493) );
  AOI32X1 U384 ( .A0(n239), .A1(n358), .A2(n557), .B0(v33), .B1(n359), .Y(n357) );
  OAI21XL U385 ( .A0(n551), .A1(n239), .B0(n4), .Y(n359) );
  XNOR2X1 U386 ( .A(n174), .B(n65), .Y(n239) );
  INVX1 U387 ( .A(n67), .Y(n65) );
  XOR2X1 U388 ( .A(n43), .B(n175), .Y(n67) );
  XNOR2X1 U389 ( .A(n519), .B(n112), .Y(n43) );
  INVX1 U390 ( .A(v25), .Y(n354) );
  OAI21XL U391 ( .A0(n6), .A1(n358), .B0(n360), .Y(n494) );
  AOI32X1 U392 ( .A0(n361), .A1(n362), .A2(n557), .B0(v41), .B1(n363), .Y(n360) );
  INVX1 U393 ( .A(v33), .Y(n358) );
  OAI222XL U394 ( .A0(v49), .A1(n97), .B0(n364), .B1(n365), .C0(n532), .C1(
        n362), .Y(n495) );
  INVX1 U395 ( .A(v41), .Y(n362) );
  AOI221X1 U396 ( .A0(n94), .A1(n78), .B0(n96), .B1(n76), .C0(n540), .Y(n364)
         );
  AOI22X1 U397 ( .A0(n76), .A1(n94), .B0(n78), .B1(n522), .Y(n97) );
  INVX1 U399 ( .A(n76), .Y(n78) );
  INVX1 U401 ( .A(n320), .Y(n318) );
  XOR2X1 U402 ( .A(n332), .B(n366), .Y(n76) );
  OAI21XL U403 ( .A0(n534), .A1(n365), .B0(n367), .Y(n496) );
  AOI32X1 U404 ( .A0(n88), .A1(n368), .A2(n557), .B0(v57), .B1(n90), .Y(n367)
         );
  OAI21XL U405 ( .A0(n551), .A1(n88), .B0(n544), .Y(n90) );
  XNOR2X1 U406 ( .A(n130), .B(n114), .Y(n88) );
  INVX1 U407 ( .A(n150), .Y(n130) );
  XNOR2X1 U408 ( .A(n295), .B(n366), .Y(n150) );
  INVX1 U409 ( .A(v49), .Y(n365) );
  OAI222XL U410 ( .A0(n79), .A1(n369), .B0(v65), .B1(n81), .C0(n532), .C1(n368), .Y(n497) );
  INVX1 U411 ( .A(v57), .Y(n368) );
  AOI22X1 U412 ( .A0(n86), .A1(n202), .B0(n85), .B1(n204), .Y(n81) );
  AOI221X1 U413 ( .A0(n86), .A1(n204), .B0(n85), .B1(n202), .C0(n540), .Y(n79)
         );
  INVX1 U420 ( .A(r2), .Y(n157) );
  OAI222XL U421 ( .A0(n370), .A1(n371), .B0(v73), .B1(n372), .C0(n532), .C1(
        n369), .Y(n498) );
  INVX1 U422 ( .A(v65), .Y(n369) );
  AOI22X1 U423 ( .A0(n521), .A1(n366), .B0(n516), .B1(n145), .Y(n372) );
  AOI221X1 U424 ( .A0(n14), .A1(n366), .B0(n12), .B1(n145), .C0(n539), .Y(n370) );
  INVX1 U426 ( .A(n145), .Y(n366) );
  OAI21XL U428 ( .A0(n6), .A1(n371), .B0(n373), .Y(n499) );
  AOI32X1 U429 ( .A0(n141), .A1(n374), .A2(n557), .B0(v81), .B1(n375), .Y(n373) );
  OAI21XL U430 ( .A0(n552), .A1(n141), .B0(n541), .Y(n375) );
  XNOR2X1 U431 ( .A(n200), .B(n145), .Y(n141) );
  INVX1 U432 ( .A(v73), .Y(n371) );
  OAI222XL U433 ( .A0(n376), .A1(n377), .B0(v89), .B1(n378), .C0(n532), .C1(
        n374), .Y(n500) );
  INVX1 U434 ( .A(v81), .Y(n374) );
  AOI22X1 U435 ( .A0(n121), .A1(n108), .B0(n287), .B1(n200), .Y(n378) );
  AOI221X1 U436 ( .A0(n287), .A1(n108), .B0(n121), .B1(n200), .C0(n537), .Y(
        n376) );
  OAI21XL U438 ( .A0(n6), .A1(n377), .B0(n379), .Y(n501) );
  AOI32X1 U439 ( .A0(n361), .A1(n380), .A2(n557), .B0(v97), .B1(n363), .Y(n379) );
  OAI21XL U440 ( .A0(n551), .A1(n361), .B0(n543), .Y(n363) );
  INVX1 U441 ( .A(v97), .Y(n380) );
  XNOR2X1 U442 ( .A(n325), .B(n50), .Y(n361) );
  XNOR2X1 U443 ( .A(n55), .B(n30), .Y(n50) );
  INVX1 U444 ( .A(n29), .Y(n30) );
  XNOR2X1 U445 ( .A(n309), .B(n174), .Y(n325) );
  INVX1 U446 ( .A(n234), .Y(n174) );
  XOR2X1 U447 ( .A(n332), .B(n200), .Y(n234) );
  INVX1 U448 ( .A(n108), .Y(n200) );
  INVX1 U450 ( .A(r7), .Y(n206) );
  XNOR2X1 U451 ( .A(message[3]), .B(n99), .Y(n332) );
  INVX1 U452 ( .A(r3), .Y(n99) );
  XNOR2X1 U453 ( .A(n320), .B(n294), .Y(n309) );
  INVX1 U454 ( .A(n295), .Y(n294) );
  XNOR2X1 U455 ( .A(message[5]), .B(n5), .Y(n295) );
  INVX1 U456 ( .A(r5), .Y(n5) );
  XNOR2X1 U457 ( .A(message[4]), .B(n313), .Y(n320) );
  INVX1 U458 ( .A(r4), .Y(n313) );
  INVX1 U459 ( .A(v89), .Y(n377) );
  INVX1 U460 ( .A(n381), .Y(n502) );
  AOI222X1 U461 ( .A0(n344), .A1(n287), .B0(n55), .B1(n121), .C0(n535), .C1(
        v97), .Y(n381) );
  NAND2X1 U465 ( .A(n555), .B(n175), .Y(n119) );
  XOR2X1 U466 ( .A(n29), .B(n145), .Y(n175) );
  INVX1 U468 ( .A(r0), .Y(n132) );
  XNOR2X1 U469 ( .A(message[1]), .B(n346), .Y(n29) );
  INVX1 U470 ( .A(r1), .Y(n346) );
  INVX1 U472 ( .A(n55), .Y(n344) );
  INVX1 U474 ( .A(r6), .Y(n244) );
  OAI22X1 U475 ( .A0(n524), .A1(n382), .B0(n548), .B1(n205), .Y(n503) );
  INVX1 U476 ( .A(message[0]), .Y(n205) );
  OAI22X1 U477 ( .A0(n524), .A1(n383), .B0(n548), .B1(n243), .Y(n504) );
  INVX1 U478 ( .A(message[1]), .Y(n243) );
  OAI22X1 U479 ( .A0(n524), .A1(n384), .B0(n548), .B1(n3), .Y(n505) );
  INVX1 U480 ( .A(message[2]), .Y(n3) );
  OAI22X1 U481 ( .A0(n524), .A1(n385), .B0(n548), .B1(n312), .Y(n506) );
  INVX1 U482 ( .A(message[3]), .Y(n312) );
  OAI22X1 U483 ( .A0(n524), .A1(n386), .B0(n548), .B1(n98), .Y(n507) );
  INVX1 U484 ( .A(message[4]), .Y(n98) );
  OAI22X1 U485 ( .A0(n524), .A1(n387), .B0(n548), .B1(n156), .Y(n508) );
  INVX1 U486 ( .A(message[5]), .Y(n156) );
  OAI22X1 U487 ( .A0(n524), .A1(n388), .B0(n548), .B1(n345), .Y(n509) );
  INVX1 U488 ( .A(message[6]), .Y(n345) );
  OAI22X1 U489 ( .A0(n524), .A1(n389), .B0(n548), .B1(n131), .Y(n510) );
  INVX1 U490 ( .A(message[7]), .Y(n131) );
  NAND2X1 U491 ( .A(n541), .B(n550), .Y(n6) );
  NAND2X1 U493 ( .A(start), .B(n390), .Y(n4) );
  OAI22X1 U494 ( .A0(sel), .A1(n133), .B0(n390), .B1(n389), .Y(code_o[7]) );
  INVX1 U495 ( .A(message_r[7]), .Y(n389) );
  INVX1 U496 ( .A(parity[7]), .Y(n133) );
  OAI22X1 U497 ( .A0(sel), .A1(n347), .B0(n390), .B1(n388), .Y(code_o[6]) );
  INVX1 U498 ( .A(message_r[6]), .Y(n388) );
  INVX1 U499 ( .A(parity[6]), .Y(n347) );
  OAI22X1 U500 ( .A0(sel), .A1(n158), .B0(n390), .B1(n387), .Y(code_o[5]) );
  INVX1 U501 ( .A(message_r[5]), .Y(n387) );
  INVX1 U502 ( .A(parity[5]), .Y(n158) );
  OAI22X1 U503 ( .A0(sel), .A1(n100), .B0(n390), .B1(n386), .Y(code_o[4]) );
  INVX1 U504 ( .A(message_r[4]), .Y(n386) );
  INVX1 U505 ( .A(parity[4]), .Y(n100) );
  OAI22X1 U506 ( .A0(sel), .A1(n314), .B0(n390), .B1(n385), .Y(code_o[3]) );
  INVX1 U507 ( .A(message_r[3]), .Y(n385) );
  INVX1 U508 ( .A(parity[3]), .Y(n314) );
  OAI22X1 U509 ( .A0(sel), .A1(n7), .B0(n390), .B1(n384), .Y(code_o[2]) );
  INVX1 U510 ( .A(message_r[2]), .Y(n384) );
  INVX1 U511 ( .A(parity[2]), .Y(n7) );
  OAI22X1 U512 ( .A0(sel), .A1(n245), .B0(n390), .B1(n383), .Y(code_o[1]) );
  INVX1 U513 ( .A(message_r[1]), .Y(n383) );
  INVX1 U514 ( .A(parity[1]), .Y(n245) );
  OAI22X1 U515 ( .A0(sel), .A1(n207), .B0(n390), .B1(n382), .Y(code_o[0]) );
  INVX1 U516 ( .A(message_r[0]), .Y(n382) );
  INVX1 U518 ( .A(parity[0]), .Y(n207) );
  DFFRHQX1 \message_r_reg[7]  ( .D(n510), .CK(clk), .RN(n569), .Q(message_r[7]) );
  DFFRHQX1 \message_r_reg[6]  ( .D(n509), .CK(clk), .RN(n569), .Q(message_r[6]) );
  DFFRHQX1 \message_r_reg[5]  ( .D(n508), .CK(clk), .RN(n569), .Q(message_r[5]) );
  DFFRHQX1 \message_r_reg[4]  ( .D(n507), .CK(clk), .RN(n569), .Q(message_r[4]) );
  DFFRHQX1 \message_r_reg[3]  ( .D(n506), .CK(clk), .RN(n569), .Q(message_r[3]) );
  DFFRHQX1 \message_r_reg[2]  ( .D(n505), .CK(clk), .RN(n569), .Q(message_r[2]) );
  DFFRHQX1 \message_r_reg[1]  ( .D(n504), .CK(clk), .RN(n569), .Q(message_r[1]) );
  DFFRHQX1 \message_r_reg[0]  ( .D(n503), .CK(clk), .RN(n569), .Q(message_r[0]) );
  DFFRHQX1 r21_reg ( .D(n468), .CK(clk), .RN(n565), .Q(v21) );
  DFFRHQX1 r25_reg ( .D(n493), .CK(clk), .RN(n568), .Q(v25) );
  DFFRHQX1 \parity_reg[6]  ( .D(n489), .CK(clk), .RN(n567), .Q(parity[6]) );
  DFFRHQX1 r44_reg ( .D(n483), .CK(clk), .RN(n567), .Q(v44) );
  DFFRHQX1 \parity_reg[3]  ( .D(n477), .CK(clk), .RN(n566), .Q(parity[3]) );
  DFFRHQX1 r85_reg ( .D(n476), .CK(clk), .RN(n566), .Q(v85) );
  DFFRHQX1 \parity_reg[1]  ( .D(n454), .CK(clk), .RN(n564), .Q(parity[1]) );
  DFFRHQX1 r15_reg ( .D(n444), .CK(clk), .RN(n563), .Q(v15) );
  DFFRHQX1 \parity_reg[0]  ( .D(n442), .CK(clk), .RN(n563), .Q(parity[0]) );
  DFFRHQX1 \parity_reg[5]  ( .D(n428), .CK(clk), .RN(n561), .Q(parity[5]) );
  DFFRHQX1 \parity_reg[7]  ( .D(n421), .CK(clk), .RN(n561), .Q(parity[7]) );
  DFFRHQX1 r101_reg ( .D(n419), .CK(clk), .RN(n560), .Q(v101) );
  DFFRHQX1 \parity_reg[4]  ( .D(n412), .CK(clk), .RN(n560), .Q(parity[4]) );
  DFFRHQX1 \parity_reg[2]  ( .D(n391), .CK(clk), .RN(n558), .Q(parity[2]) );
  DFFRHQX1 r89_reg ( .D(n501), .CK(clk), .RN(n569), .Q(v89) );
  DFFRHQX1 r73_reg ( .D(n499), .CK(clk), .RN(n568), .Q(v73) );
  DFFRHQX1 r65_reg ( .D(n498), .CK(clk), .RN(n568), .Q(v65) );
  DFFRHQX1 r84_reg ( .D(n488), .CK(clk), .RN(n567), .Q(v84) );
  DFFRHQX1 r76_reg ( .D(n487), .CK(clk), .RN(n567), .Q(v76) );
  DFFRHQX1 r68_reg ( .D(n486), .CK(clk), .RN(n567), .Q(v68) );
  DFFRHQX1 r60_reg ( .D(n485), .CK(clk), .RN(n567), .Q(v60) );
  DFFRHQX1 r52_reg ( .D(n484), .CK(clk), .RN(n567), .Q(v52) );
  DFFRHQX1 r36_reg ( .D(n482), .CK(clk), .RN(n567), .Q(v36) );
  DFFRHQX1 r28_reg ( .D(n481), .CK(clk), .RN(n567), .Q(v28) );
  DFFRHQX1 r20_reg ( .D(n480), .CK(clk), .RN(n566), .Q(v20) );
  DFFRHQX1 r77_reg ( .D(n475), .CK(clk), .RN(n566), .Q(v77) );
  DFFRHQX1 r61_reg ( .D(n473), .CK(clk), .RN(n566), .Q(v61) );
  DFFRHQX1 r45_reg ( .D(n471), .CK(clk), .RN(n566), .Q(v45) );
  DFFRHQX1 r37_reg ( .D(n470), .CK(clk), .RN(n565), .Q(v37) );
  DFFRHQX1 r86_reg ( .D(n465), .CK(clk), .RN(n565), .Q(v86) );
  DFFRHQX1 r78_reg ( .D(n464), .CK(clk), .RN(n565), .Q(v78) );
  DFFRHQX1 r62_reg ( .D(n462), .CK(clk), .RN(n565), .Q(v62) );
  DFFRHQX1 r30_reg ( .D(n458), .CK(clk), .RN(n564), .Q(v30) );
  DFFRHQX1 r14_reg ( .D(n456), .CK(clk), .RN(n564), .Q(v14) );
  DFFRHQX1 r87_reg ( .D(n453), .CK(clk), .RN(n564), .Q(v87) );
  DFFRHQX1 r79_reg ( .D(n452), .CK(clk), .RN(n564), .Q(v79) );
  DFFRHQX1 r71_reg ( .D(n451), .CK(clk), .RN(n564), .Q(v71) );
  DFFRHQX1 r47_reg ( .D(n448), .CK(clk), .RN(n563), .Q(v47) );
  DFFRHQX1 r31_reg ( .D(n446), .CK(clk), .RN(n563), .Q(v31) );
  DFFRHQX1 r74_reg ( .D(n438), .CK(clk), .RN(n562), .Q(v74) );
  DFFRHQX1 r66_reg ( .D(n437), .CK(clk), .RN(n562), .Q(v66) );
  DFFRHQX1 r58_reg ( .D(n436), .CK(clk), .RN(n562), .Q(v58) );
  DFFRHQX1 r26_reg ( .D(n432), .CK(clk), .RN(n562), .Q(v26) );
  DFFRHQX1 r18_reg ( .D(n431), .CK(clk), .RN(n562), .Q(v18) );
  DFFRHQX1 r24_reg ( .D(n425), .CK(clk), .RN(n561), .Q(v24) );
  DFFRHQX1 r8_reg ( .D(n423), .CK(clk), .RN(n561), .Q(v8) );
  DFFRHQX1 r93_reg ( .D(n418), .CK(clk), .RN(n560), .Q(v93) );
  DFFRHQX1 r27_reg ( .D(n416), .CK(clk), .RN(n560), .Q(v27) );
  DFFRHQX1 r99_reg ( .D(n411), .CK(clk), .RN(n560), .Q(v99) );
  DFFRHQX1 r83_reg ( .D(n409), .CK(clk), .RN(n559), .Q(v83) );
  DFFRHQX1 r75_reg ( .D(n408), .CK(clk), .RN(n559), .Q(v75) );
  DFFRHQX1 r67_reg ( .D(n407), .CK(clk), .RN(n559), .Q(v67) );
  DFFRHQX1 r80_reg ( .D(n402), .CK(clk), .RN(n559), .Q(v80) );
  DFFRHQX1 r64_reg ( .D(n400), .CK(clk), .RN(n558), .Q(v64) );
  DFFRHQX1 r94_reg ( .D(n394), .CK(clk), .RN(n558), .Q(v94) );
  DFFRHQX1 r100_reg ( .D(n393), .CK(clk), .RN(n558), .Q(v100) );
  DFFRHQX1 r92_reg ( .D(n392), .CK(clk), .RN(n558), .Q(v92) );
  DFFRHQX1 r49_reg ( .D(n496), .CK(clk), .RN(n568), .Q(v49) );
  DFFRHQX1 r51_reg ( .D(n405), .CK(clk), .RN(n559), .Q(v51) );
  DFFRHQX1 r81_reg ( .D(n500), .CK(clk), .RN(n568), .Q(v81) );
  DFFRHQX1 r57_reg ( .D(n497), .CK(clk), .RN(n568), .Q(v57) );
  DFFRHQX1 r41_reg ( .D(n495), .CK(clk), .RN(n568), .Q(v41) );
  DFFRHQX1 r33_reg ( .D(n494), .CK(clk), .RN(n568), .Q(v33) );
  DFFRHQX1 r29_reg ( .D(n469), .CK(clk), .RN(n565), .Q(v29) );
  DFFRHQX1 r54_reg ( .D(n461), .CK(clk), .RN(n565), .Q(v54) );
  DFFRHQX1 r46_reg ( .D(n460), .CK(clk), .RN(n564), .Q(v46) );
  DFFRHQX1 r22_reg ( .D(n457), .CK(clk), .RN(n564), .Q(v22) );
  DFFRHQX1 r63_reg ( .D(n450), .CK(clk), .RN(n563), .Q(v63) );
  DFFRHQX1 r55_reg ( .D(n449), .CK(clk), .RN(n563), .Q(v55) );
  DFFRHQX1 r23_reg ( .D(n445), .CK(clk), .RN(n563), .Q(v23) );
  DFFRHQX1 r90_reg ( .D(n440), .CK(clk), .RN(n562), .Q(v90) );
  DFFRHQX1 r50_reg ( .D(n435), .CK(clk), .RN(n562), .Q(v50) );
  DFFRHQX1 r42_reg ( .D(n434), .CK(clk), .RN(n562), .Q(v42) );
  DFFRHQX1 r34_reg ( .D(n433), .CK(clk), .RN(n562), .Q(v34) );
  DFFRHQX1 r19_reg ( .D(n415), .CK(clk), .RN(n560), .Q(v19) );
  DFFRHQX1 r91_reg ( .D(n410), .CK(clk), .RN(n559), .Q(v91) );
  DFFRHQX1 r59_reg ( .D(n406), .CK(clk), .RN(n559), .Q(v59) );
  DFFRHQX1 r72_reg ( .D(n401), .CK(clk), .RN(n559), .Q(v72) );
  DFFRHQX1 r56_reg ( .D(n399), .CK(clk), .RN(n558), .Q(v56) );
  DFFRHQX1 r48_reg ( .D(n398), .CK(clk), .RN(n558), .Q(v48) );
  DFFRHQX1 r102_reg ( .D(n395), .CK(clk), .RN(n558), .Q(v102) );
  DFFRHQX1 r17_reg ( .D(n492), .CK(clk), .RN(n568), .Q(v17) );
  DFFRHQX1 r9_reg ( .D(n491), .CK(clk), .RN(n568), .Q(v9) );
  DFFRHQX1 r12_reg ( .D(n479), .CK(clk), .RN(n566), .Q(v12) );
  DFFRHQX1 r69_reg ( .D(n474), .CK(clk), .RN(n566), .Q(v69) );
  DFFRHQX1 r13_reg ( .D(n467), .CK(clk), .RN(n565), .Q(v13) );
  DFFRHQX1 r70_reg ( .D(n463), .CK(clk), .RN(n565), .Q(v70) );
  DFFRHQX1 r38_reg ( .D(n459), .CK(clk), .RN(n564), .Q(v38) );
  DFFRHQX1 r39_reg ( .D(n447), .CK(clk), .RN(n563), .Q(v39) );
  DFFRHQX1 r82_reg ( .D(n439), .CK(clk), .RN(n562), .Q(v82) );
  DFFRHQX1 r10_reg ( .D(n430), .CK(clk), .RN(n561), .Q(v10) );
  DFFRHQX1 r40_reg ( .D(n427), .CK(clk), .RN(n561), .Q(v40) );
  DFFRHQX1 r32_reg ( .D(n426), .CK(clk), .RN(n561), .Q(v32) );
  DFFRHQX1 r16_reg ( .D(n424), .CK(clk), .RN(n561), .Q(v16) );
  DFFRHQX1 r96_reg ( .D(n420), .CK(clk), .RN(n560), .Q(v96) );
  DFFRHQX1 r88_reg ( .D(n417), .CK(clk), .RN(n560), .Q(v88) );
  DFFRHQX1 r11_reg ( .D(n414), .CK(clk), .RN(n560), .Q(v11) );
  DFFRHQX1 r43_reg ( .D(n404), .CK(clk), .RN(n559), .Q(v43) );
  DFFRHQX1 r95_reg ( .D(n396), .CK(clk), .RN(n558), .Q(v95) );
  DFFRHQX1 r53_reg ( .D(n472), .CK(clk), .RN(n566), .Q(v53) );
  DFFRHQX1 r35_reg ( .D(n403), .CK(clk), .RN(n559), .Q(v35) );
  DFFRHQX1 r103_reg ( .D(n397), .CK(clk), .RN(n558), .Q(v103) );
  DFFRHQX1 r97_reg ( .D(n502), .CK(clk), .RN(n569), .Q(v97) );
  DFFRHQX1 r98_reg ( .D(n441), .CK(clk), .RN(n563), .Q(v98) );
  DFFRHQX1 r4_reg ( .D(n478), .CK(clk), .RN(n566), .Q(r4) );
  DFFRHQX1 r5_reg ( .D(n466), .CK(clk), .RN(n565), .Q(r5) );
  DFFRHQX1 r7_reg ( .D(n443), .CK(clk), .RN(n563), .Q(r7) );
  DFFRHQX1 r3_reg ( .D(n413), .CK(clk), .RN(n560), .Q(r3) );
  DFFRHQX1 r1_reg ( .D(n490), .CK(clk), .RN(n567), .Q(r1) );
  DFFRHQX1 r6_reg ( .D(n455), .CK(clk), .RN(n564), .Q(r6) );
  DFFRHQX1 r2_reg ( .D(n429), .CK(clk), .RN(n561), .Q(r2) );
  DFFRHQX1 r0_reg ( .D(n422), .CK(clk), .RN(n561), .Q(r0) );
  INVX1 U519 ( .A(n515), .Y(n511) );
  INVX1 U520 ( .A(n513), .Y(n512) );
  BUFX3 U521 ( .A(n114), .Y(n513) );
  INVX1 U522 ( .A(n249), .Y(n514) );
  BUFX3 U523 ( .A(n86), .Y(n515) );
  BUFX3 U524 ( .A(n14), .Y(n516) );
  INVX1 U525 ( .A(n118), .Y(n517) );
  BUFX3 U526 ( .A(n94), .Y(n518) );
  INVX1 U527 ( .A(n344), .Y(n519) );
  INVX1 U528 ( .A(n116), .Y(n520) );
  INVX1 U529 ( .A(n296), .Y(n521) );
  BUFX3 U530 ( .A(n96), .Y(n522) );
  INVX1 U531 ( .A(n535), .Y(n524) );
  INVX1 U532 ( .A(n535), .Y(n525) );
  INVX1 U533 ( .A(n535), .Y(n526) );
  INVX1 U534 ( .A(n536), .Y(n527) );
  INVX1 U535 ( .A(n536), .Y(n528) );
  INVX1 U536 ( .A(n536), .Y(n529) );
  INVX1 U537 ( .A(n536), .Y(n531) );
  INVX1 U538 ( .A(n536), .Y(n530) );
  INVX1 U539 ( .A(n535), .Y(n532) );
  INVX1 U540 ( .A(n536), .Y(n533) );
  INVX1 U541 ( .A(n535), .Y(n534) );
  NOR2X1 U542 ( .A(n174), .B(n549), .Y(n14) );
  NOR2X1 U543 ( .A(n549), .B(n301), .Y(n75) );
  INVX1 U544 ( .A(n119), .Y(n287) );
  INVX1 U545 ( .A(n556), .Y(n549) );
  INVX1 U546 ( .A(n556), .Y(n548) );
  INVX1 U547 ( .A(n555), .Y(n550) );
  INVX1 U548 ( .A(n542), .Y(n537) );
  INVX1 U549 ( .A(n6), .Y(n535) );
  INVX1 U550 ( .A(n555), .Y(n551) );
  INVX1 U551 ( .A(n555), .Y(n552) );
  INVX1 U552 ( .A(n6), .Y(n536) );
  INVX1 U553 ( .A(n556), .Y(n554) );
  INVX1 U554 ( .A(n523), .Y(n553) );
  NOR2X1 U555 ( .A(n548), .B(n234), .Y(n12) );
  XNOR2X1 U556 ( .A(n43), .B(n234), .Y(n228) );
  NOR2X1 U557 ( .A(n549), .B(n318), .Y(n94) );
  NOR2X1 U558 ( .A(n548), .B(n294), .Y(n66) );
  NOR2X1 U559 ( .A(n309), .B(n550), .Y(n77) );
  NOR2X1 U560 ( .A(n175), .B(n549), .Y(n121) );
  NOR2X1 U561 ( .A(n549), .B(n30), .Y(n204) );
  INVX1 U562 ( .A(n85), .Y(n86) );
  INVX1 U563 ( .A(n541), .Y(n538) );
  INVX1 U564 ( .A(n541), .Y(n539) );
  INVX1 U565 ( .A(n541), .Y(n540) );
  INVX1 U566 ( .A(n547), .Y(n555) );
  INVX1 U567 ( .A(n547), .Y(n556) );
  INVX1 U568 ( .A(n546), .Y(n542) );
  INVX1 U569 ( .A(n546), .Y(n545) );
  INVX1 U570 ( .A(n546), .Y(n543) );
  INVX1 U571 ( .A(n546), .Y(n544) );
  INVX1 U572 ( .A(n547), .Y(n557) );
  INVX1 U573 ( .A(n114), .Y(n112) );
  XOR2X1 U574 ( .A(n332), .B(n112), .Y(n85) );
  NOR2X1 U575 ( .A(n320), .B(n549), .Y(n96) );
  NOR2X1 U576 ( .A(n295), .B(n550), .Y(n64) );
  NOR2X1 U577 ( .A(n29), .B(n549), .Y(n202) );
  XOR2X1 U578 ( .A(n332), .B(n344), .Y(n242) );
  INVX1 U579 ( .A(n546), .Y(n541) );
  INVX1 U580 ( .A(n4), .Y(n546) );
  INVX1 U581 ( .A(n523), .Y(n547) );
  INVX1 U582 ( .A(n571), .Y(n558) );
  INVX1 U583 ( .A(n571), .Y(n559) );
  INVX1 U584 ( .A(n571), .Y(n560) );
  INVX1 U585 ( .A(n570), .Y(n561) );
  INVX1 U586 ( .A(n570), .Y(n562) );
  INVX1 U587 ( .A(n570), .Y(n563) );
  INVX1 U588 ( .A(n570), .Y(n564) );
  INVX1 U589 ( .A(n571), .Y(n565) );
  INVX1 U590 ( .A(n570), .Y(n566) );
  INVX1 U591 ( .A(n571), .Y(n567) );
  INVX1 U592 ( .A(n570), .Y(n568) );
  INVX1 U593 ( .A(n571), .Y(n569) );
  XNOR2X1 U594 ( .A(message[6]), .B(n244), .Y(n55) );
  XNOR2X1 U595 ( .A(message[0]), .B(n132), .Y(n145) );
  XNOR2X1 U596 ( .A(message[2]), .B(n157), .Y(n114) );
  XNOR2X1 U597 ( .A(message[7]), .B(n206), .Y(n108) );
  INVX1 U598 ( .A(sel), .Y(n390) );
  AND2X2 U599 ( .A(sel), .B(start), .Y(n523) );
  INVX1 U600 ( .A(reset), .Y(n571) );
  INVX1 U601 ( .A(reset), .Y(n570) );
endmodule

