module multiplier_column2_p16(b,P1,P2,P3,P4,P5,P6,P7,P8,
                                P9,P10,P11,P12,P13,P14,P15,P16);

input [12:0]b;
output [12:0]P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16; 

//wire[415:0]P;

wire	[207:0]P;

wire BBM1,BBM2,BBM3,BBM4,BBM5,BBM6,BBM7,BBM8,BBM9,BBM10,
BBM11,BBM12,BBM13,BBM14,BBM15,BBM16,BBM17,BBM18,BBM19,BBM20,
BBM21,BBM22,BBM23,BBM24,BBM25,BBM26,BBM27,BBM28,BBM29,BBM30,
BBM31,BBM32,BBM33,BBM34,BBM35,BBM36,BBM37,BBM38,BBM39,BBM40,
BBM41,BBM42,BBM43,BBM44,BBM45,BBM46,BBM47,BBM48,BBM49,BBM50,
BBM51,BBM52,BBM53,BBM54,BBM55,BBM56,BBM57,BBM58,BBM59,BBM60,
BBM61,BBM62,BBM63,BBM64,BBM65,BBM66,BBM67,BBM68,BBM69,BBM70,
BBM71,BBM72,BBM73,BBM74,BBM75,BBM76,BBM77,BBM78,BBM79,BBM80,
BBM81,BBM82,BBM83,BBM84,BBM85,BBM86,BBM87,BBM88,BBM89,BBM90,
BBM91,BBM92,BBM93,BBM94,BBM95,BBM96,BBM97,BBM98,BBM99,BBM100,
BBM101,BBM102,BBM103,BBM104,BBM105,BBM106,BBM107,BBM108,BBM109,BBM110,
BBM111,BBM112,BBM113,BBM114,BBM115,BBM116,BBM117,BBM118,BBM119,BBM120,
BBM121,BBM122,BBM123,BBM124,BBM125,BBM126,BBM127,BBM128,BBM129,BBM130,
BBM131,BBM132,BBM133,BBM134,BBM135,BBM136,BBM137,BBM138,BBM139,BBM140,
BBM141,BBM142,BBM143,BBM144,BBM145,BBM146,BBM147,BBM148,BBM149,BBM150,
BBM151,BBM152,BBM153,BBM154,BBM155,BBM156,BBM157,BBM158,BBM159,BBM160,
BBM161,BBM162,BBM163,BBM164,BBM165,BBM166,BBM167,BBM168,BBM169,BBM170,
BBM171,BBM172,BBM173,BBM174,BBM175,BBM176,BBM177,BBM178,BBM179,BBM180,
BBM181,BBM182,BBM183,BBM184,BBM185,BBM186,BBM187,BBM188,BBM189,BBM190,
BBM191,BBM192,BBM193,BBM194,BBM195,BBM196,BBM197,BBM198,BBM199,BBM200,
BBM201,BBM202,BBM203,BBM204,BBM205,BBM206,BBM207,BBM208;


assign BBM1=BBM8^BBM142;
assign BBM2=BBM19^BBM171^b[8];
assign BBM3=BBM16^BBM143;
assign BBM5=BBM45^BBM144;
assign BBM6=BBM29^BBM176;
assign BBM8=BBM49^BBM177;
assign BBM9=BBM29^b[6];
assign BBM10=BBM47^BBM177;
assign BBM16=BBM34^b[6];
assign BBM17=BBM75^b[0]^b[6];
assign BBM18=BBM76^b[3]^b[11];
assign BBM19=BBM49^b[7];
assign BBM20=BBM76^BBM179;
assign BBM21=BBM83^BBM145;
assign BBM29=BBM57^BBM178;
assign BBM34=BBM113^b[1]^b[4];
assign BBM35=BBM74^b[1];
assign BBM36=BBM75^b[1];
assign BBM37=BBM96^b[3]^b[4];
assign BBM40=BBM115^BBM180;
assign BBM43=BBM106^b[0]^b[1];
assign BBM45=BBM114^BBM168;
assign BBM46=BBM146^BBM147;
assign BBM47=BBM73^b[10];
assign BBM49=BBM113^b[0]^b[5];
assign BBM53=BBM117^b[3];
assign BBM54=BBM138^BBM162;
assign BBM55=BBM146^BBM184;
assign BBM57=BBM139^BBM181;
assign BBM58=BBM114^b[0];
assign BBM60=BBM141^BBM168;
assign BBM64=BBM129^b[3]^b[5];
assign BBM67=BBM116^b[10];
assign BBM71=BBM144^b[5]^b[10];
assign BBM72=BBM116^b[7];
assign BBM73=BBM117^b[5];
assign BBM74=BBM115^b[5];
assign BBM75=BBM140^BBM183;
assign BBM76=BBM100^b[1];
assign BBM82=BBM154^BBM157;
assign BBM83=BBM158^BBM159;
assign BBM84=BBM129^b[8];
assign BBM85=BBM160^BBM162;
assign BBM86=BBM131^b[6];
assign BBM88=BBM145^b[12];
assign BBM89=BBM133^b[4];
assign BBM96=BBM155^b[0]^b[9];
assign BBM100=BBM131^b[12];
assign BBM101=BBM143^b[1];
assign BBM104=BBM178^b[6]^b[10];
assign BBM105=BBM167^BBM168;
assign BBM106=BBM175^b[7]^b[12];
assign BBM113=BBM153^BBM184;
assign BBM114=BBM142^b[12];
assign BBM115=BBM137^b[4];
assign BBM116=BBM160^BBM173;
assign BBM117=BBM147^b[4];
assign BBM128=BBM153^b[2];
assign BBM129=BBM153^b[9];
assign BBM130=BBM155^b[10];
assign BBM131=BBM157^b[7];
assign BBM133=BBM159^b[5];
assign BBM137=BBM183^b[12];
assign BBM138=BBM165^b[11];
assign BBM139=BBM170^b[8];
assign BBM140=BBM160^b[11];
assign BBM141=BBM181^b[4];
assign BBM143=BBM177^b[7];
assign BBM144=BBM166^b[4];
assign BBM145=BBM162^b[3];
assign BBM146=BBM172^b[0];
assign BBM147=BBM163^b[12];
assign BBM4=b[0]^b[2]^b[3]^b[4]^b[5]^b[7]^b[8]^b[10]^b[11]^b[12];
assign BBM7=b[1]^b[3]^b[4]^b[5]^b[6]^b[8]^b[9]^b[11]^b[12];
assign BBM11=b[0]^b[4]^b[6]^b[7]^b[8]^b[9]^b[11]^b[12];
assign BBM12=b[2]^b[4]^b[5]^b[6]^b[7]^b[9]^b[10]^b[12];
assign BBM13=b[0]^b[4]^b[6]^b[7]^b[8]^b[9]^b[11]^b[12];
assign BBM14=b[2]^b[4]^b[5]^b[6]^b[7]^b[9]^b[10]^b[12];
assign BBM15=b[0]^b[4]^b[6]^b[7]^b[8]^b[9]^b[11]^b[12];
assign BBM22=b[0]^b[2]^b[6]^b[8]^b[9]^b[10]^b[11];
assign BBM23=b[1]^b[3]^b[7]^b[9]^b[10]^b[11]^b[12];
assign BBM24=b[1]^b[5]^b[7]^b[8]^b[9]^b[10]^b[12];
assign BBM25=b[1]^b[3]^b[7]^b[9]^b[10]^b[11]^b[12];
assign BBM26=b[3]^b[5]^b[6]^b[7]^b[8]^b[10]^b[11];
assign BBM27=b[0]^b[2]^b[6]^b[8]^b[9]^b[10]^b[11];
assign BBM28=b[1]^b[5]^b[7]^b[8]^b[9]^b[10]^b[12];
assign BBM30=b[3]^b[5]^b[6]^b[7]^b[8]^b[10]^b[11];
assign BBM31=b[0]^b[2]^b[6]^b[8]^b[9]^b[10]^b[11];
assign BBM32=b[1]^b[3]^b[7]^b[9]^b[10]^b[11]^b[12];
assign BBM33=b[1]^b[5]^b[7]^b[8]^b[9]^b[10]^b[12];
assign BBM38=b[1]^b[2]^b[4]^b[5]^b[10]^b[12];
assign BBM39=b[0]^b[1]^b[3]^b[4]^b[9]^b[11];
assign BBM41=b[1]^b[2]^b[4]^b[5]^b[10]^b[12];
assign BBM42=b[0]^b[1]^b[3]^b[4]^b[9]^b[11];
assign BBM44=b[2]^b[4]^b[8]^b[10]^b[11]^b[12];
assign BBM48=b[2]^b[4]^b[8]^b[10]^b[11]^b[12];
assign BBM50=b[1]^b[2]^b[4]^b[5]^b[10]^b[12];
assign BBM51=b[0]^b[1]^b[3]^b[4]^b[9]^b[11];
assign BBM52=b[2]^b[4]^b[8]^b[10]^b[11]^b[12];
assign BBM56=b[3]^b[4]^b[6]^b[7]^b[12];
assign BBM59=b[2]^b[3]^b[5]^b[6]^b[11];
assign BBM61=b[0]^b[2]^b[3]^b[8]^b[10];
assign BBM62=b[3]^b[4]^b[6]^b[7]^b[12];
assign BBM63=b[2]^b[3]^b[5]^b[6]^b[11];
assign BBM65=b[0]^b[1]^b[6]^b[8]^b[12];
assign BBM66=b[0]^b[2]^b[3]^b[8]^b[10];
assign BBM68=b[3]^b[5]^b[9]^b[11]^b[12];
assign BBM69=b[0]^b[1]^b[6]^b[8]^b[12];
assign BBM70=b[3]^b[5]^b[9]^b[11]^b[12];
assign BBM77=b[3]^b[4]^b[6]^b[7]^b[12];
assign BBM78=b[2]^b[3]^b[5]^b[6]^b[11];
assign BBM79=b[0]^b[2]^b[3]^b[8]^b[10];
assign BBM80=b[0]^b[1]^b[6]^b[8]^b[12];
assign BBM81=b[3]^b[5]^b[9]^b[11]^b[12];
assign BBM87=b[0]^b[9]^b[10]^b[12];
assign BBM90=b[7]^b[8]^b[10]^b[11];
assign BBM91=b[8]^b[9]^b[11]^b[12];
assign BBM92=b[5]^b[6]^b[8]^b[9];
assign BBM93=b[6]^b[7]^b[9]^b[10];
assign BBM94=b[0]^b[9]^b[10]^b[12];
assign BBM95=b[8]^b[9]^b[11]^b[12];
assign BBM97=b[4]^b[5]^b[7]^b[8];
assign BBM98=b[7]^b[8]^b[10]^b[11];
assign BBM99=b[6]^b[7]^b[9]^b[10];
assign BBM102=b[5]^b[6]^b[8]^b[9];
assign BBM103=b[4]^b[5]^b[7]^b[8];
assign BBM107=b[1]^b[2]^b[7]^b[9];
assign BBM108=b[4]^b[6]^b[10]^b[12];
assign BBM109=b[0]^b[5]^b[7]^b[11];
assign BBM110=b[1]^b[2]^b[7]^b[9];
assign BBM111=b[0]^b[5]^b[7]^b[11];
assign BBM112=b[4]^b[6]^b[10]^b[12];
assign BBM118=b[7]^b[8]^b[10]^b[11];
assign BBM119=b[0]^b[9]^b[10]^b[12];
assign BBM120=b[8]^b[9]^b[11]^b[12];
assign BBM121=b[5]^b[6]^b[8]^b[9];
assign BBM122=b[6]^b[7]^b[9]^b[10];
assign BBM123=b[4]^b[5]^b[7]^b[8];
assign BBM124=b[7]^b[8]^b[10]^b[11];
assign BBM125=b[1]^b[2]^b[7]^b[9];
assign BBM126=b[4]^b[6]^b[10]^b[12];
assign BBM127=b[0]^b[5]^b[7]^b[11];
assign BBM132=b[2]^b[11]^b[12];
assign BBM134=b[1]^b[10]^b[11];
assign BBM135=b[2]^b[11]^b[12];
assign BBM136=b[1]^b[10]^b[11];
assign BBM142=b[1]^b[6]^b[8];
assign BBM148=b[9]^b[11]^b[12];
assign BBM149=b[7]^b[9]^b[10];
assign BBM150=b[5]^b[7]^b[8];
assign BBM151=b[2]^b[11]^b[12];
assign BBM152=b[1]^b[10]^b[11];
assign BBM153=b[11]^b[12];
assign BBM154=b[0]^b[12];
assign BBM155=b[1]^b[11];
assign BBM156=b[3]^b[12];
assign BBM157=b[9]^b[10];
assign BBM158=b[10]^b[11];
assign BBM159=b[7]^b[8];
assign BBM160=b[8]^b[9];
assign BBM161=b[3]^b[12];
assign BBM162=b[5]^b[6];
assign BBM163=b[6]^b[7];
assign BBM164=b[3]^b[12];
assign BBM165=b[2]^b[3];
assign BBM166=b[3]^b[9];
assign BBM167=b[0]^b[7];
assign BBM168=b[5]^b[11];
assign BBM169=b[6]^b[11];
assign BBM170=b[0]^b[11];
assign BBM171=b[2]^b[4];
assign BBM172=b[2]^b[8];
assign BBM173=b[1]^b[3];
assign BBM174=b[3]^b[6];
assign BBM175=b[2]^b[5];
assign BBM176=b[1]^b[10];
assign BBM177=b[2]^b[9];
assign BBM178=b[4]^b[12];
assign BBM179=b[5]^b[8];
assign BBM180=b[8]^b[11];
assign BBM181=b[7]^b[9];
assign BBM182=b[5]^b[11];
assign BBM183=b[2]^b[10];
assign BBM184=b[3]^b[10];
assign BBM185=b[7]^b[9];
assign BBM186=b[11]^b[12];
assign BBM187=b[7]^b[8];
assign BBM188=b[11]^b[12];
assign BBM189=b[3]^b[12];
assign BBM190=b[3]^b[12];
assign BBM191=b[5]^b[11];
assign BBM192=b[7]^b[9];
assign BBM193=b[11];

assign P[1]=BBM153;
assign P[2]=BBM154;
assign P[3]=BBM155;
assign P[4]=BBM128;
assign P[5]=BBM156;
assign P[14]=BBM157;
assign P[15]=BBM158;
assign P[16]=BBM129;
assign P[17]=BBM82;
assign P[18]=BBM130;
assign P[19]=BBM128;
assign P[20]=BBM156;
assign P[27]=BBM159;
assign P[28]=BBM160;
assign P[29]=BBM131;
assign P[30]=BBM83;
assign P[31]=BBM84;
assign P[32]=BBM82;
assign P[33]=BBM130;
assign P[34]=BBM128;
assign P[35]=BBM156;
assign P[40]=BBM162;
assign P[41]=BBM163;
assign P[42]=BBM133;
assign P[43]=BBM85;
assign P[44]=BBM86;
assign P[45]=BBM83;
assign P[46]=BBM84;
assign P[47]=BBM82;
assign P[48]=BBM130;
assign P[49]=BBM128;
assign P[50]=BBM156;
assign P[52]=BBM156;
assign P[53]=BBM156^b[4];
assign P[55]=BBM88;
assign P[56]=BBM53;
assign P[57]=BBM89;
assign P[58]=BBM85;
assign P[59]=BBM86;
assign P[60]=BBM83;
assign P[61]=BBM84;
assign P[62]=BBM82;
assign P[63]=BBM130;
assign P[64]=BBM128;
assign P[65]=BBM130;
assign P[66]=BBM137^b[1];
assign P[67]=BBM138;
assign P[68]=BBM34;
assign P[69]=BBM35;
assign P[70]=BBM54;
assign P[71]=BBM53;
assign P[72]=BBM89;
assign P[73]=BBM85;
assign P[74]=BBM86;
assign P[75]=BBM83;
assign P[76]=BBM84;
assign P[77]=BBM82;
assign P[78]=BBM84;
assign P[79]=BBM139^b[10];
assign P[80]=BBM96^b[12];
assign P[81]=BBM36;
assign P[82]=BBM55;
assign P[83]=BBM37;
assign P[84]=BBM35;
assign P[85]=BBM54;
assign P[86]=BBM53;
assign P[87]=BBM89;
assign P[88]=BBM85;
assign P[89]=BBM86;
assign P[90]=BBM83;
assign P[91]=BBM86;
assign P[92]=BBM140^b[6];
assign P[93]=BBM100;
assign P[94]=BBM57^b[6];
assign P[95]=BBM58;
assign P[96]=BBM101;
assign P[97]=BBM55;
assign P[98]=BBM37;
assign P[99]=BBM35;
assign P[100]=BBM54;
assign P[101]=BBM53;
assign P[102]=BBM89;
assign P[103]=BBM85;
assign P[104]=BBM89;
assign P[105]=BBM141^b[6];
assign P[106]=BBM133^b[10];
assign P[107]=BBM60^b[6];
assign P[108]=BBM104;
assign P[109]=BBM105;
assign P[110]=BBM58;
assign P[111]=BBM101;
assign P[112]=BBM55;
assign P[113]=BBM37;
assign P[114]=BBM35;
assign P[115]=BBM54;
assign P[116]=BBM53;
assign P[117]=BBM54;
assign P[118]=BBM106^b[4]^b[11];
assign P[119]=BBM88^b[8];
assign P[120]=BBM60^BBM165;
assign P[121]=BBM40;
assign P[122]=BBM64;
assign P[123]=BBM104;
assign P[124]=BBM105;
assign P[125]=BBM58;
assign P[126]=BBM101;
assign P[127]=BBM55;
assign P[128]=BBM37;
assign P[129]=BBM35;
assign P[130]=BBM37;
assign P[131]=BBM8;
assign P[132]=BBM16;
assign P[133]=BBM43^BBM166;
assign P[134]=BBM17;
assign P[135]=BBM18;
assign P[136]=BBM40;
assign P[137]=BBM64;
assign P[138]=BBM104;
assign P[139]=BBM105;
assign P[140]=BBM58;
assign P[141]=BBM101;
assign P[142]=BBM55;
assign P[143]=BBM101;
assign P[144]=BBM67^BBM167;
assign P[145]=BBM36^b[4];
assign P[146]=BBM19^b[1];
assign P[147]=BBM9;
assign P[148]=BBM20;
assign P[149]=BBM17;
assign P[150]=BBM18;
assign P[151]=BBM40;
assign P[152]=BBM64;
assign P[153]=BBM104;
assign P[154]=BBM105;
assign P[155]=BBM58;
assign P[156]=BBM105;
assign P[157]=BBM45^b[7];
assign P[158]=BBM46^b[9];
assign P[159]=BBM67^BBM168;
assign P[160]=BBM10;
assign P[161]=BBM21;
assign P[162]=BBM9;
assign P[163]=BBM20;
assign P[164]=BBM17;
assign P[165]=BBM18;
assign P[166]=BBM40;
assign P[167]=BBM64;
assign P[168]=BBM104;
assign P[169]=BBM64;
assign P[170]=BBM71^BBM169;
assign P[171]=BBM47^BBM170;
assign P[172]=BBM72^b[6];
assign P[173]=BBM2;
assign P[174]=BBM5;
assign P[175]=BBM10;
assign P[176]=BBM21;
assign P[177]=BBM9;
assign P[178]=BBM20;
assign P[179]=BBM17;
assign P[180]=BBM18;
assign P[181]=BBM40;
assign P[182]=BBM18;
assign P[183]=BBM72^BBM171;
assign P[184]=BBM71^BBM172;
assign P[185]=BBM73^b[1];
assign P[186]=BBM1;
assign P[187]=BBM3;
assign P[188]=BBM2;
assign P[189]=BBM5;
assign P[190]=BBM10;
assign P[191]=BBM21;
assign P[192]=BBM9;
assign P[193]=BBM20;
assign P[194]=BBM17;
assign P[195]=BBM20;
assign P[196]=BBM43^BBM169;
assign P[197]=BBM46^BBM173;
assign P[198]=BBM74^b[3];
assign P[199]=BBM6^BBM174;
assign P[200]=BBM6^BBM175;
assign P[201]=BBM1;
assign P[202]=BBM3;
assign P[203]=BBM2;
assign P[204]=BBM5;
assign P[205]=BBM10;
assign P[206]=BBM21;
assign P[207]=BBM9;
assign P[0]=b[11];
assign P[6]=b[4];
assign P[7]=b[5];
assign P[8]=b[6];
assign P[9]=b[7];
assign P[10]=b[8];
assign P[11]=b[9];
assign P[12]=b[10];
assign P[13]=b[9];
assign P[21]=b[4];
assign P[22]=b[5];
assign P[23]=b[6];
assign P[24]=b[7];
assign P[25]=b[8];
assign P[26]=b[7];
assign P[36]=b[4];
assign P[37]=b[5];
assign P[38]=b[6];
assign P[39]=b[5];
assign P[51]=b[4];
assign P[54]=b[4]^b[5];


assign P1[12:0]=P[12:0];
assign P2[12:0]=P[25:13];
assign P3[12:0]=P[38:26];
assign P4[12:0]=P[51:39];
assign P5[12:0]=P[64:52];
assign P6[12:0]=P[77:65];
assign P7[12:0]=P[90:78];
assign P8[12:0]=P[103:91];
assign P9[12:0]=P[116:104];
assign P10[12:0]=P[129:117];
assign P11[12:0]=P[142:130];
assign P12[12:0]=P[155:143];
assign P13[12:0]=P[168:156];
assign P14[12:0]=P[181:169];
assign P15[12:0]=P[194:182];
assign P16[12:0]=P[207:195];








endmodule
