module multiplier(a,b,c);

input [12:0]a,b;
output [12:0]c;

wire [12:0]c,d;
wire [11:0]e;

 //-----d=Lb------------------------------

assign d[0]=(a[0]&b[0]);
assign d[1]=(a[1]&b[0])^(a[0]&b[1]);
assign d[2]=(a[2]&b[0])^(a[1]&b[1])^(a[0]&b[2]);
assign d[3]=(a[3]&b[0])^(a[2]&b[1])^(a[1]&b[2])^(a[0]&b[3]);
assign d[4]=(a[4]&b[0])^(a[3]&b[1])^(a[2]&b[2])^(a[1]&b[3])^(a[0]&b[4]);
assign d[5]=(a[5]&b[0])^(a[4]&b[1])^(a[3]&b[2])^(a[2]&b[3])^(a[1]&b[4])^(a[0]&b[5]);
assign d[6]=(a[6]&b[0])^(a[5]&b[1])^(a[4]&b[2])^(a[3]&b[3])^(a[2]&b[4])^(a[1]&b[5])^(a[0]&b[6]);
assign d[7]=(a[7]&b[0])^(a[6]&b[1])^(a[5]&b[2])^(a[4]&b[3])^(a[3]&b[4])^(a[2]&b[5])^(a[1]&b[6])^(a[0]&b[7]);
assign d[8]=(a[8]&b[0])^(a[7]&b[1])^(a[6]&b[2])^(a[5]&b[3])^(a[4]&b[4])^(a[3]&b[5])^(a[2]&b[6])^(a[1]&b[7])^(a[0]&b[8]);
assign d[9]=(a[9]&b[0])^(a[8]&b[1])^(a[7]&b[2])^(a[6]&b[3])^(a[5]&b[4])^(a[4]&b[5])^(a[3]&b[6])^(a[2]&b[7])^(a[1]&b[8])^(a[0]&b[9]);
assign d[10]=(a[10]&b[0])^(a[9]&b[1])^(a[8]&b[2])^(a[7]&b[3])^(a[6]&b[4])^(a[5]&b[5])^(a[4]&b[6])^(a[3]&b[7])^(a[2]&b[8])^(a[1]&b[9])^(a[0]&b[10]);
assign d[11]=(a[11]&b[0])^(a[10]&b[1])^(a[9]&b[2])^(a[8]&b[3])^(a[7]&b[4])^(a[6]&b[5])^(a[5]&b[6])^(a[4]&b[7])^(a[3]&b[8])^(a[2]&b[9])^(a[1]&b[10])^(a[0]&b[11]);
assign d[12]=(a[12]&b[0])^(a[11]&b[1])^(a[10]&b[2])^(a[9]&b[3])^(a[8]&b[4])^(a[7]&b[5])^(a[6]&b[6])^(a[5]&b[7])^(a[4]&b[8])^(a[3]&b[9])^(a[2]&b[10])^(a[1]&b[11])^(a[0]&b[12]);




//--------e=Ub----------------------------------------
assign e[0]=(a[12]&b[1])^(a[11]&b[2])^(a[10]&b[3])^(a[9]&b[4])^(a[8]&b[5])^(a[7]&b[6])^(a[6]&b[7])^(a[5]&b[8])^(a[4]&b[9])^(a[3]&b[10])^(a[2]&b[11])^(a[1]&b[12]);
assign e[1]=(a[12]&b[2])^(a[11]&b[3])^(a[10]&b[4])^(a[9]&b[5])^(a[8]&b[6])^(a[7]&b[7])^(a[6]&b[8])^(a[5]&b[9])^(a[4]&b[10])^(a[3]&b[11])^(a[2]&b[12]);
assign e[2]=(a[12]&b[3])^(a[11]&b[4])^(a[10]&b[5])^(a[9]&b[6])^(a[8]&b[7])^(a[7]&b[8])^(a[6]&b[9])^(a[5]&b[10])^(a[4]&b[11])^(a[3]&b[12]);
assign e[3]=(a[12]&b[4])^(a[11]&b[5])^(a[10]&b[6])^(a[9]&b[7])^(a[8]&b[8])^(a[7]&b[9])^(a[6]&b[10])^(a[5]&b[11])^(a[4]&b[12]);
assign e[4]=(a[12]&b[5])^(a[11]&b[6])^(a[10]&b[7])^(a[9]&b[8])^(a[8]&b[9])^(a[7]&b[10])^(a[6]&b[11])^(a[5]&b[12]);
assign e[5]=(a[12]&b[6])^(a[11]&b[7])^(a[10]&b[8])^(a[9]&b[9])^(a[8]&b[10])^(a[7]&b[11])^(a[6]&b[12]);
assign e[6]=(a[12]&b[7])^(a[11]&b[8])^(a[10]&b[9])^(a[9]&b[10])^(a[8]&b[11])^(a[7]&b[12]);
assign e[7]=(a[12]&b[8])^(a[11]&b[9])^(a[10]&b[10])^(a[9]&b[11])^(a[8]&b[12]);
assign e[8]=(a[12]&b[9])^(a[11]&b[10])^(a[10]&b[11])^(a[9]&b[12]);
assign e[9]=(a[12]&b[10])^(a[11]&b[11])^(a[10]&b[12]);
assign e[10]=(a[12]&b[11])^(a[11]&b[12]);
assign e[11]=(a[12]&b[12]);

//----------c=d+Q^t+e--------------------------------------
assign c[0]=d[0]^e[0] ^e[9] ^e[10] ;
assign c[1]=d[1]^e[0] ^e[1] ^e[9] ^e[11] ;
assign c[2]=d[2]^e[1] ^e[2] ^e[10] ;
assign c[3]=d[3]^e[0] ^e[2] ^e[3] ^e[9] ^e[10] ^e[11] ;
assign c[4]=d[4]^e[0] ^e[1] ^e[3] ^e[4] ^e[9] ^e[11] ;
assign c[5]=d[5]^e[1] ^e[2] ^e[4] ^e[5] ^e[10] ;
assign c[6]=d[6]^e[2] ^e[3] ^e[5] ^e[6] ^e[11] ;
assign c[7]=d[7]^e[3] ^e[4] ^e[6] ^e[7] ;
assign c[8]=d[8]^e[4] ^e[5] ^e[7] ^e[8] ;
assign c[9]=d[9]^e[5] ^e[6] ^e[8] ^e[9] ;
assign c[10]=d[10]^e[6] ^e[7] ^e[9] ^e[10] ;
assign c[11]=d[11]^e[7] ^e[8] ^e[10] ^e[11] ;
assign c[12]=d[12]^e[8] ^e[9] ^e[11] ;



  

endmodule
