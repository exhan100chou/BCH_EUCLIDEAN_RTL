module multiplier_column6_p16(b,P1,P2,P3,P4,P5,P6,P7,P8,
                                P9,P10,P11,P12,P13,P14,P15,P16);

input [12:0]b;
output [12:0]P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16; 

//wire[415:0]P;

wire	[207:0]P;

wire BBM1,BBM2,BBM3,BBM4,BBM5,BBM6,BBM7,BBM8,BBM9,BBM10,
BBM11,BBM12,BBM13,BBM14,BBM15,BBM16,BBM17,BBM18,BBM19,BBM20,
BBM21,BBM22,BBM23,BBM24,BBM25,BBM26,BBM27,BBM28,BBM29,BBM30,
BBM31,BBM32,BBM33,BBM34,BBM35,BBM36,BBM37,BBM38,BBM39,BBM40,
BBM41,BBM42,BBM43,BBM44,BBM45,BBM46,BBM47,BBM48,BBM49,BBM50,
BBM51,BBM52,BBM53,BBM54,BBM55,BBM56,BBM57,BBM58,BBM59,BBM60,
BBM61,BBM62,BBM63,BBM64,BBM65,BBM66,BBM67,BBM68,BBM69,BBM70,
BBM71,BBM72,BBM73,BBM74,BBM75,BBM76,BBM77,BBM78,BBM79,BBM80,
BBM81,BBM82,BBM83,BBM84,BBM85,BBM86,BBM87,BBM88,BBM89,BBM90,
BBM91,BBM92,BBM93,BBM94,BBM95,BBM96,BBM97,BBM98,BBM99,BBM100,
BBM101,BBM102,BBM103,BBM104,BBM105,BBM106,BBM107,BBM108,BBM109,BBM110,
BBM111,BBM112,BBM113,BBM114,BBM115,BBM116,BBM117,BBM118,BBM119,BBM120,
BBM121,BBM122,BBM123,BBM124,BBM125,BBM126,BBM127,BBM128,BBM129,BBM130,
BBM131,BBM132,BBM133,BBM134,BBM135,BBM136,BBM137,BBM138,BBM139,BBM140,
BBM141,BBM142,BBM143,BBM144,BBM145,BBM146,BBM147,BBM148,BBM149,BBM150,
BBM151,BBM152,BBM153,BBM154,BBM155,BBM156,BBM157,BBM158,BBM159,BBM160,
BBM161,BBM162,BBM163,BBM164,BBM165,BBM166,BBM167,BBM168,BBM169,BBM170,
BBM171,BBM172,BBM173,BBM174,BBM175,BBM176,BBM177,BBM178,BBM179,BBM180,
BBM181,BBM182,BBM183,BBM184,BBM185,BBM186,BBM187,BBM188,BBM189,BBM190,
BBM191,BBM192,BBM193,BBM194,BBM195,BBM196,BBM197,BBM198,BBM199,BBM200,
BBM201,BBM202,BBM203,BBM204,BBM205,BBM206,BBM207,BBM208,BBM209,BBM210,
BBM211,BBM212,BBM213,BBM214,BBM215,BBM216,BBM217,BBM218;

assign BBM1=BBM9^BBM184;
assign BBM2=BBM16^BBM182^b[6];
assign BBM3=BBM13^b[0]^b[7];
assign BBM4=BBM9^b[7];
assign BBM5=BBM24^BBM185;
assign BBM6=BBM27^BBM186;
assign BBM7=BBM27^BBM187;
assign BBM8=BBM26^b[1]^b[4];
assign BBM9=BBM15^b[3]^b[5];
assign BBM10=BBM39^BBM177;
assign BBM11=BBM45^BBM188;
assign BBM12=BBM46^b[5]^b[11];
assign BBM13=BBM31^b[3]^b[5];
assign BBM14=BBM40^b[8];
assign BBM15=BBM47^b[6];
assign BBM16=BBM48^BBM183;
assign BBM17=BBM62^BBM189;
assign BBM18=BBM47^b[5];
assign BBM19=BBM46^b[9];
assign BBM20=BBM57^BBM179;
assign BBM21=BBM45^b[9];
assign BBM22=BBM64^BBM191;
assign BBM23=BBM80^BBM192;
assign BBM24=BBM72^BBM193;
assign BBM25=BBM61^BBM185;
assign BBM26=BBM65^BBM194;
assign BBM27=BBM81^BBM195;
assign BBM28=BBM59^b[10];
assign BBM29=BBM108^BBM194;
assign BBM30=BBM95^BBM185;
assign BBM31=BBM106^BBM182;
assign BBM32=BBM99^BBM193;
assign BBM33=BBM82^b[2];
assign BBM34=BBM108^b[0]^b[2];
assign BBM35=BBM88^BBM195;
assign BBM36=BBM109^BBM197;
assign BBM37=BBM81^b[11];
assign BBM38=BBM68^b[8];
assign BBM39=BBM110^BBM188;
assign BBM40=BBM98^BBM198;
assign BBM41=BBM82^b[4];
assign BBM42=BBM109^BBM199;
assign BBM43=BBM83^b[11];
assign BBM44=BBM83^b[8];
assign BBM45=BBM80^b[8];
assign BBM46=BBM105^BBM200;
assign BBM47=BBM94^b[9]^b[11];
assign BBM48=BBM125^BBM165;
assign BBM49=BBM96^b[11];
assign BBM50=BBM107^b[7];
assign BBM51=BBM111^b[5];
assign BBM52=BBM112^b[6];
assign BBM53=BBM143^b[0]^b[9];
assign BBM54=BBM113^b[4];
assign BBM55=BBM144^BBM201;
assign BBM56=BBM120^b[2];
assign BBM57=BBM101^b[5];
assign BBM58=BBM126^BBM194;
assign BBM59=BBM114^b[5];
assign BBM60=BBM144^b[4]^b[8];
assign BBM61=BBM115^b[11];
assign BBM62=BBM91^b[9];
assign BBM63=BBM90^b[3];
assign BBM64=BBM117^b[7];
assign BBM65=BBM86^b[0];
assign BBM67=BBM113^b[5];
assign BBM68=BBM146^BBM201;
assign BBM69=BBM119^b[12];
assign BBM70=BBM120^b[0];
assign BBM71=BBM103^b[1];
assign BBM72=BBM111^b[1];
assign BBM73=BBM119^b[9];
assign BBM74=BBM120^b[10];
assign BBM75=BBM117^b[5];
assign BBM76=BBM115^b[2];
assign BBM77=BBM119^b[1];
assign BBM79=BBM88^b[4];
assign BBM80=BBM133^BBM189;
assign BBM81=BBM89^b[1];
assign BBM82=BBM112^b[7];
assign BBM83=BBM135^b[6]^b[7];
assign BBM85=BBM137^b[11];
assign BBM86=BBM138^b[12];
assign BBM87=BBM139^b[0];
assign BBM88=BBM135^b[10];
assign BBM89=BBM136^b[8];
assign BBM90=BBM124^b[6];
assign BBM91=BBM130^b[4];
assign BBM92=BBM131^b[5];
assign BBM93=BBM149^b[7];
assign BBM94=BBM174^BBM200;
assign BBM95=BBM125^b[0];
assign BBM96=BBM171^BBM172;
assign BBM97=BBM151^b[12];
assign BBM98=BBM168^BBM202;
assign BBM99=BBM132^b[11];
assign BBM100=BBM152^b[11];
assign BBM101=BBM153^b[1];
assign BBM102=BBM154^b[5];
assign BBM103=BBM151^b[10];
assign BBM104=BBM140^b[0];
assign BBM105=BBM176^BBM180;
assign BBM106=BBM147^b[12];
assign BBM107=BBM153^b[3];
assign BBM108=BBM155^b[1];
assign BBM109=BBM152^b[10];
assign BBM110=BBM138^b[0];
assign BBM111=BBM188^b[9]^b[11];
assign BBM112=BBM169^b[0]^b[12];
assign BBM113=BBM149^b[8];
assign BBM114=BBM135^b[4];
assign BBM115=BBM154^b[7];
assign BBM117=BBM134^b[4];
assign BBM119=BBM145^b[8];
assign BBM120=BBM155^b[4];
assign BBM124=BBM183^b[10];
assign BBM125=BBM166^b[1];
assign BBM126=BBM179^b[11];
assign BBM127=BBM170^b[5];
assign BBM128=BBM183^b[6];
assign BBM129=BBM168^b[8];
assign BBM130=BBM192^b[6];
assign BBM131=BBM173^b[7];
assign BBM132=BBM168^b[6];
assign BBM133=BBM181^b[3];
assign BBM134=BBM166^b[0];
assign BBM135=BBM176^b[12];
assign BBM136=BBM197^b[5];
assign BBM137=BBM162^b[10];
assign BBM138=BBM163^b[11];
assign BBM139=BBM192^b[9];
assign BBM140=BBM164^b[1];
assign BBM143=BBM191^b[11];
assign BBM144=BBM164^b[3];
assign BBM145=BBM167^b[2];
assign BBM146=BBM178^b[6];
assign BBM147=BBM166^b[8];
assign BBM149=BBM176^b[9];
assign BBM150=BBM173^b[1];
assign BBM151=BBM201^b[4];
assign BBM152=BBM171^b[0];
assign BBM153=BBM188^b[12];
assign BBM154=BBM208^b[6];
assign BBM155=BBM163^b[3];
assign BBM66=b[2]^b[3]^b[7]^b[10]^b[11];
assign BBM78=b[2]^b[3]^b[4]^b[8]^b[9];
assign BBM84=b[2]^b[3]^b[4]^b[8]^b[9];
assign BBM116=b[4]^b[6]^b[10]^b[12];
assign BBM118=b[8]^b[9]^b[11]^b[12];
assign BBM121=b[2]^b[3]^b[7]^b[8];
assign BBM122=b[4]^b[5]^b[7]^b[8];
assign BBM123=b[3]^b[4]^b[8]^b[9];
assign BBM141=b[5]^b[6]^b[8];
assign BBM142=b[6]^b[7]^b[9];
assign BBM148=b[1]^b[2]^b[12];
assign BBM156=b[0]^b[10]^b[11];
assign BBM157=b[8]^b[9]^b[11];
assign BBM158=b[2]^b[3]^b[7];
assign BBM159=b[4]^b[5]^b[7];
assign BBM160=b[6]^b[7]^b[9];
assign BBM161=b[1]^b[2]^b[12];
assign BBM162=b[7]^b[8];
assign BBM163=b[8]^b[9];
assign BBM164=b[11]^b[12];
assign BBM165=b[3]^b[12];
assign BBM166=b[10]^b[11];
assign BBM167=b[3]^b[7];
assign BBM168=b[5]^b[10];
assign BBM169=b[1]^b[8];
assign BBM170=b[6]^b[8];
assign BBM171=b[3]^b[6];
assign BBM172=b[2]^b[5];
assign BBM173=b[0]^b[11];
assign BBM174=b[2]^b[8];
assign BBM175=b[8]^b[11];
assign BBM176=b[1]^b[2];
assign BBM177=b[7]^b[12];
assign BBM178=b[2]^b[12];
assign BBM179=b[2]^b[3];
assign BBM180=b[3]^b[4];
assign BBM181=b[0]^b[5];
assign BBM182=b[2]^b[4];
assign BBM183=b[7]^b[9];
assign BBM184=b[1]^b[12];
assign BBM185=b[5]^b[12];
assign BBM186=b[0]^b[3];
assign BBM187=b[2]^b[10];
assign BBM188=b[4]^b[6];
assign BBM189=b[2]^b[7];
assign BBM190=b[2]^b[3];
assign BBM191=b[1]^b[3];
assign BBM192=b[10]^b[12];
assign BBM193=b[3]^b[8];
assign BBM194=b[7]^b[10];
assign BBM195=b[6]^b[9];
assign BBM196=b[5]^b[12];
assign BBM197=b[4]^b[7];
assign BBM198=b[9]^b[12];
assign BBM199=b[2]^b[9];
assign BBM200=b[0]^b[10];
assign BBM201=b[5]^b[9];
assign BBM202=b[1]^b[7];
assign BBM203=b[3]^b[6];
assign BBM204=b[4]^b[9];
assign BBM205=b[7]^b[9];
assign BBM206=b[10]^b[11];
assign BBM207=b[5]^b[10];
assign BBM208=b[0]^b[1];
assign BBM209=b[4]^b[6];
assign BBM210=b[10]^b[11];
assign BBM211=b[8]^b[9];
assign BBM212=b[1]^b[2];
assign BBM213=b[5]^b[10];
assign BBM214=b[3]^b[6];
assign BBM215=b[2]^b[3];
assign BBM216=b[7]^b[9];
assign BBM217=b[10]^b[11];
assign BBM218=b[7];
assign P[1]=BBM162;
assign P[2]=BBM163;
assign P[3]=BBM124;
assign P[4]=BBM85;
assign P[5]=BBM86;
assign P[6]=BBM87;
assign P[7]=BBM125;
assign P[8]=BBM164^b[2];
assign P[9]=BBM165;
assign P[13]=BBM125;
assign P[14]=BBM88;
assign P[15]=BBM126;
assign P[16]=BBM48^b[4];
assign P[17]=BBM28;
assign P[18]=BBM49;
assign P[19]=BBM50;
assign P[20]=BBM89;
assign P[21]=BBM127^b[9];
assign P[22]=BBM90;
assign P[23]=BBM85;
assign P[24]=BBM86;
assign P[25]=BBM87;
assign P[26]=BBM89;
assign P[27]=BBM128^b[4];
assign P[28]=BBM129^b[7];
assign P[29]=BBM51^b[7];
assign P[30]=BBM91;
assign P[31]=BBM92;
assign P[32]=BBM52;
assign P[33]=BBM93;
assign P[34]=BBM94^b[3];
assign P[35]=BBM53^b[4];
assign P[36]=BBM28;
assign P[37]=BBM49;
assign P[38]=BBM50;
assign P[39]=BBM93;
assign P[40]=BBM29^b[0];
assign P[41]=BBM54^BBM166;
assign P[42]=BBM30^BBM167;
assign P[43]=BBM10;
assign P[44]=BBM14;
assign P[45]=BBM15;
assign P[46]=BBM16;
assign P[47]=BBM31;
assign P[48]=BBM55;
assign P[49]=BBM91;
assign P[50]=BBM92;
assign P[51]=BBM52;
assign P[52]=BBM16;
assign P[53]=BBM54^BBM167;
assign P[54]=BBM56^BBM168;
assign P[55]=BBM57^b[7];
assign P[56]=BBM1;
assign P[57]=BBM2;
assign P[58]=BBM3;
assign P[59]=BBM5;
assign P[60]=BBM17^b[5];
assign P[61]=BBM32^b[7];
assign P[62]=BBM10;
assign P[63]=BBM14;
assign P[64]=BBM15;
assign P[65]=BBM5;
assign P[66]=BBM58^BBM169;
assign P[67]=BBM56^BBM164;
assign P[68]=BBM95^BBM170;
assign P[69]=BBM11;
assign P[70]=BBM6;
assign P[71]=BBM7;
assign P[72]=BBM4;
assign P[73]=BBM8^BBM171;
assign P[74]=BBM8^BBM172;
assign P[75]=BBM1;
assign P[76]=BBM2;
assign P[77]=BBM3;
assign P[78]=BBM4;
assign P[79]=BBM59;
assign P[80]=BBM96;
assign P[81]=BBM18^b[4];
assign P[82]=BBM33;
assign P[83]=BBM34;
assign P[84]=BBM19;
assign P[85]=BBM12;
assign P[86]=BBM20^BBM173;
assign P[87]=BBM20^b[7];
assign P[88]=BBM11;
assign P[89]=BBM6;
assign P[90]=BBM7;
assign P[91]=BBM12;
assign P[92]=BBM130;
assign P[93]=BBM131;
assign P[94]=BBM13;
assign P[95]=BBM35;
assign P[96]=BBM58;
assign P[97]=BBM60;
assign P[98]=BBM97;
assign P[99]=BBM132^b[0];
assign P[100]=BBM61;
assign P[101]=BBM33;
assign P[102]=BBM34;
assign P[103]=BBM19;
assign P[104]=BBM97;
assign P[105]=BBM62^b[0];
assign P[106]=BBM98^b[11];
assign P[107]=BBM51^BBM174;
assign P[108]=BBM36;
assign P[109]=BBM37;
assign P[110]=BBM38;
assign P[111]=BBM63;
assign P[112]=BBM64^b[8];
assign P[113]=BBM65^b[1]^b[5];
assign P[114]=BBM35;
assign P[115]=BBM58;
assign P[116]=BBM60;
assign P[117]=BBM63;
assign P[118]=BBM39^b[3];
assign P[119]=BBM40^b[4];
assign P[120]=BBM21^b[11];
assign P[121]=BBM41;
assign P[122]=BBM67;
assign P[123]=BBM42;
assign P[124]=BBM22;
assign P[125]=BBM59^BBM175;
assign P[126]=BBM68^b[3];
assign P[127]=BBM36;
assign P[128]=BBM37;
assign P[129]=BBM38;
assign P[130]=BBM22;
assign P[131]=BBM23^b[8];
assign P[132]=BBM24;
assign P[133]=BBM55^BBM176;
assign P[134]=BBM43;
assign P[135]=BBM69;
assign P[136]=BBM70;
assign P[137]=BBM71;
assign P[138]=BBM99^b[2];
assign P[139]=BBM100^BBM177;
assign P[140]=BBM41;
assign P[141]=BBM67;
assign P[142]=BBM42;
assign P[143]=BBM71;
assign P[144]=BBM72^b[2];
assign P[145]=BBM23;
assign P[146]=BBM32^b[9];
assign P[147]=BBM25;
assign P[148]=BBM44;
assign P[149]=BBM73;
assign P[150]=BBM74;
assign P[151]=BBM75^b[9];
assign P[152]=BBM30^b[6];
assign P[153]=BBM43;
assign P[154]=BBM69;
assign P[155]=BBM70;
assign P[156]=BBM74;
assign P[157]=BBM133^BBM175;
assign P[158]=BBM101^b[9];
assign P[159]=BBM21^b[4];
assign P[160]=BBM102;
assign P[161]=BBM76;
assign P[162]=BBM77;
assign P[163]=BBM56;
assign P[164]=BBM103^b[3];
assign P[165]=BBM75^b[6];
assign P[166]=BBM25;
assign P[167]=BBM44;
assign P[168]=BBM73;
assign P[169]=BBM56;
assign P[170]=BBM129^b[2];
assign P[171]=BBM100^b[9];
assign P[172]=BBM29^BBM178;
assign P[173]=BBM134;
assign P[174]=BBM104;
assign P[175]=BBM135;
assign P[176]=BBM179;
assign P[177]=BBM180;
assign P[178]=BBM181^b[4];
assign P[179]=BBM102;
assign P[180]=BBM76;
assign P[181]=BBM77;
assign P[182]=BBM179;
assign P[183]=BBM182;
assign P[184]=BBM133;
assign P[185]=BBM105^b[6];
assign P[186]=BBM136;
assign P[187]=BBM127;
assign P[188]=BBM128;
assign P[189]=BBM137;
assign P[190]=BBM138;
assign P[191]=BBM139;
assign P[192]=BBM134;
assign P[193]=BBM104;
assign P[194]=BBM135;
assign P[195]=BBM137;
assign P[196]=BBM124^b[11];
assign P[197]=BBM106;
assign P[198]=BBM26;
assign P[199]=BBM140^BBM183;
assign P[200]=BBM94^b[12];
assign P[201]=BBM53;
assign P[202]=BBM79;
assign P[203]=BBM126^b[5];
assign P[204]=BBM107;
assign P[205]=BBM136;
assign P[206]=BBM127;
assign P[207]=BBM128;
assign P[0]=b[7];
assign P[10]=b[4];
assign P[11]=b[5];
assign P[12]=b[6];



assign P1[12:0]=P[12:0];
assign P2[12:0]=P[25:13];
assign P3[12:0]=P[38:26];
assign P4[12:0]=P[51:39];
assign P5[12:0]=P[64:52];
assign P6[12:0]=P[77:65];
assign P7[12:0]=P[90:78];
assign P8[12:0]=P[103:91];
assign P9[12:0]=P[116:104];
assign P10[12:0]=P[129:117];
assign P11[12:0]=P[142:130];
assign P12[12:0]=P[155:143];
assign P13[12:0]=P[168:156];
assign P14[12:0]=P[181:169];
assign P15[12:0]=P[194:182];
assign P16[12:0]=P[207:195];








endmodule
