module multiplier_column8_p16(b,P1,P2,P3,P4,P5,P6,P7,P8,
                                P9,P10,P11,P12,P13,P14,P15,P16);

input [12:0]b;
output [12:0]P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16; 

//wire[415:0]P;

wire	[207:0]P;

wire BBM1,BBM2,BBM3,BBM4,BBM5,BBM6,BBM7,BBM8,BBM9,BBM10,
BBM11,BBM12,BBM13,BBM14,BBM15,BBM16,BBM17,BBM18,BBM19,BBM20,
BBM21,BBM22,BBM23,BBM24,BBM25,BBM26,BBM27,BBM28,BBM29,BBM30,
BBM31,BBM32,BBM33,BBM34,BBM35,BBM36,BBM37,BBM38,BBM39,BBM40,
BBM41,BBM42,BBM43,BBM44,BBM45,BBM46,BBM47,BBM48,BBM49,BBM50,
BBM51,BBM52,BBM53,BBM54,BBM55,BBM56,BBM57,BBM58,BBM59,BBM60,
BBM61,BBM62,BBM63,BBM64,BBM65,BBM66,BBM67,BBM68,BBM69,BBM70,
BBM71,BBM72,BBM73,BBM74,BBM75,BBM76,BBM77,BBM78,BBM79,BBM80,
BBM81,BBM82,BBM83,BBM84,BBM85,BBM86,BBM87,BBM88,BBM89,BBM90,
BBM91,BBM92,BBM93,BBM94,BBM95,BBM96,BBM97,BBM98,BBM99,BBM100,
BBM101,BBM102,BBM103,BBM104,BBM105,BBM106,BBM107,BBM108,BBM109,BBM110,
BBM111,BBM112,BBM113,BBM114,BBM115,BBM116,BBM117,BBM118,BBM119,BBM120,
BBM121,BBM122,BBM123,BBM124,BBM125,BBM126,BBM127,BBM128,BBM129,BBM130,
BBM131,BBM132,BBM133,BBM134,BBM135,BBM136,BBM137,BBM138,BBM139,BBM140,
BBM141,BBM142,BBM143,BBM144,BBM145,BBM146,BBM147,BBM148,BBM149,BBM150,
BBM151,BBM152,BBM153,BBM154,BBM155,BBM156,BBM157,BBM158,BBM159,BBM160,
BBM161,BBM162,BBM163,BBM164,BBM165,BBM166,BBM167,BBM168,BBM169,BBM170,
BBM171,BBM172,BBM173,BBM174,BBM175,BBM176,BBM177,BBM178,BBM179,BBM180,
BBM181,BBM182,BBM183,BBM184,BBM185,BBM186,BBM187,BBM188,BBM189,BBM190,
BBM191,BBM192,BBM193,BBM194,BBM195,BBM196,BBM197,BBM198,BBM199,BBM200,
BBM201,BBM202,BBM203,BBM204,BBM205,BBM206,BBM207,BBM208,BBM209,BBM210,
BBM211,BBM212,BBM213,BBM214,BBM215,BBM216,BBM217,BBM218,BBM219,BBM220,
BBM221,BBM222,BBM223,BBM224,BBM225,BBM226,BBM227,BBM228,BBM229,BBM230,
BBM231;

assign BBM1=BBM4^BBM186;
assign BBM2=BBM5^BBM167;
assign BBM3=BBM24^BBM188;
assign BBM4=BBM25^BBM176;
assign BBM5=BBM42^BBM189;
assign BBM6=BBM11^b[3];
assign BBM7=BBM43^BBM190;
assign BBM8=BBM43^BBM191;
assign BBM9=BBM26^BBM181;
assign BBM10=BBM44^b[0];
assign BBM11=BBM33^b[2];
assign BBM12=BBM41^b[12];
assign BBM13=BBM48^BBM193;
assign BBM14=BBM39^b[0];
assign BBM15=BBM45^b[4];
assign BBM16=BBM46^b[2];
assign BBM17=BBM47^BBM210;
assign BBM18=BBM46^b[3];
assign BBM19=BBM44^b[2];
assign BBM20=BBM53^BBM167;
assign BBM21=BBM51^BBM190;
assign BBM22=BBM59^b[5];
assign BBM23=BBM60^b[1];
assign BBM24=BBM83^BBM194;
assign BBM25=BBM59^b[9];
assign BBM26=BBM54^b[3];
assign BBM27=BBM57^b[0];
assign BBM28=BBM58^b[3];
assign BBM29=BBM62^b[3];
assign BBM30=BBM63^b[11];
assign BBM31=BBM62^b[1];
assign BBM32=BBM84^BBM195;
assign BBM33=BBM64^b[7];
assign BBM34=BBM92^BBM183;
assign BBM35=BBM79^BBM177;
assign BBM36=BBM60^b[3];
assign BBM37=BBM63^b[1];
assign BBM38=BBM78^BBM174;
assign BBM39=BBM93^BBM197;
assign BBM40=BBM56^b[4];
assign BBM41=BBM75^b[1]^b[4];
assign BBM42=BBM88^BBM197;
assign BBM43=BBM102^BBM184^b[7];
assign BBM44=BBM98^BBM153;
assign BBM45=BBM64^b[2];
assign BBM46=BBM81^BBM179;
assign BBM47=BBM116^BBM198;
assign BBM48=BBM74^b[6];
assign BBM49=BBM69^b[5];
assign BBM50=BBM92^b[6];
assign BBM51=BBM82^b[2];
assign BBM52=BBM77^b[3];
assign BBM53=BBM123^b[0]^b[6];
assign BBM54=BBM86^b[8];
assign BBM55=BBM108^BBM199;
assign BBM56=BBM95^b[11];
assign BBM57=BBM93^b[9];
assign BBM58=BBM72^b[6];
assign BBM59=BBM123^BBM163;
assign BBM60=BBM95^b[8];
assign BBM62=BBM107^BBM172;
assign BBM63=BBM124^BBM164;
assign BBM64=BBM91^b[5];
assign BBM65=BBM134^BBM202;
assign BBM66=BBM125^b[6];
assign BBM67=BBM119^b[4];
assign BBM68=BBM120^b[5];
assign BBM69=BBM106^b[12];
assign BBM70=BBM136^b[0]^b[3];
assign BBM71=BBM126^b[2];
assign BBM72=BBM103^b[0];
assign BBM73=BBM147^BBM177;
assign BBM74=BBM113^b[12];
assign BBM75=BBM104^b[8];
assign BBM76=BBM149^BBM199;
assign BBM77=BBM135^BBM204;
assign BBM78=BBM126^b[0];
assign BBM79=BBM140^BBM194;
assign BBM80=BBM112^b[0];
assign BBM81=BBM115^b[1];
assign BBM82=BBM125^b[7];
assign BBM83=BBM152^BBM170;
assign BBM84=BBM122^b[0];
assign BBM85=BBM139^BBM198;
assign BBM86=BBM138^BBM180;
assign BBM87=BBM154^BBM207;
assign BBM88=BBM101^b[12];
assign BBM89=BBM126^b[6];
assign BBM90=BBM118^b[0];
assign BBM91=BBM117^b[6];
assign BBM92=BBM131^BBM169;
assign BBM93=BBM137^BBM173;
assign BBM95=BBM99^b[5];
assign BBM96=BBM150^b[9];
assign BBM97=BBM142^b[10];
assign BBM98=BBM143^b[12];
assign BBM99=BBM131^b[7];
assign BBM100=BBM154^b[2];
assign BBM101=BBM170^b[2]^b[8];
assign BBM102=BBM148^b[6];
assign BBM103=BBM129^b[4];
assign BBM104=BBM174^BBM197;
assign BBM105=BBM134^b[5];
assign BBM106=BBM153^b[3];
assign BBM107=BBM156^b[4];
assign BBM108=BBM161^BBM170;
assign BBM109=BBM162^BBM210;
assign BBM111=BBM177^BBM211;
assign BBM112=BBM174^b[4]^b[8];
assign BBM113=BBM158^b[7];
assign BBM115=BBM181^BBM206;
assign BBM116=BBM150^b[3];
assign BBM117=BBM160^b[12];
assign BBM118=BBM156^b[10];
assign BBM119=BBM160^b[3];
assign BBM120=BBM158^b[12];
assign BBM121=BBM165^BBM176;
assign BBM122=BBM141^b[12];
assign BBM123=BBM165^BBM218;
assign BBM124=BBM151^b[4];
assign BBM125=BBM168^BBM186;
assign BBM126=BBM182^BBM215;
assign BBM129=BBM211^b[5];
assign BBM130=BBM166^b[8];
assign BBM131=BBM171^b[10];
assign BBM132=BBM209^b[6];
assign BBM133=BBM178^b[6];
assign BBM134=BBM218^b[0];
assign BBM135=BBM171^b[5];
assign BBM136=BBM167^b[8];
assign BBM137=BBM169^b[4];
assign BBM138=BBM168^b[6];
assign BBM139=BBM206^b[0];
assign BBM140=BBM210^b[5];
assign BBM141=BBM172^b[7];
assign BBM142=BBM162^b[9];
assign BBM143=BBM194^b[9];
assign BBM144=BBM170^b[11];
assign BBM145=BBM164^b[1];
assign BBM147=BBM166^b[11];
assign BBM148=BBM172^b[11];
assign BBM149=BBM189^b[5];
assign BBM150=BBM161^b[8];
assign BBM151=BBM174^b[0];
assign BBM152=BBM204^b[9];
assign BBM153=BBM162^b[4];
assign BBM154=BBM167^b[7];
assign BBM156=BBM194^b[12];
assign BBM157=BBM166^b[9];
assign BBM158=BBM190^b[2];
assign BBM160=BBM199^b[0];
assign BBM61=b[1]^b[2]^b[6]^b[7]^b[8]^b[12];
assign BBM94=b[1]^b[4]^b[5]^b[9]^b[10];
assign BBM110=b[6]^b[7]^b[9]^b[10];
assign BBM114=b[2]^b[3]^b[7]^b[8];
assign BBM127=b[4]^b[8]^b[10]^b[11];
assign BBM128=b[7]^b[9]^b[10]^b[12];
assign BBM146=b[7]^b[8]^b[10];
assign BBM155=b[0]^b[7]^b[11];
assign BBM159=b[5]^b[6]^b[8];
assign BBM161=b[5]^b[6];
assign BBM162=b[6]^b[7];
assign BBM163=b[1]^b[10];
assign BBM164=b[2]^b[12];
assign BBM165=b[3]^b[12];
assign BBM166=b[7]^b[10];
assign BBM167=b[1]^b[9];
assign BBM168=b[1]^b[12];
assign BBM169=b[1]^b[2];
assign BBM170=b[0]^b[10];
assign BBM171=b[9]^b[12];
assign BBM172=b[2]^b[5];
assign BBM173=b[3]^b[10];
assign BBM174=b[3]^b[9];
assign BBM175=b[3]^b[4];
assign BBM176=b[4]^b[6];
assign BBM177=b[2]^b[3];
assign BBM178=b[10]^b[12];
assign BBM179=b[6]^b[8];
assign BBM180=b[2]^b[7];
assign BBM181=b[9]^b[10];
assign BBM182=b[4]^b[11];
assign BBM183=b[3]^b[8];
assign BBM184=b[0]^b[9];
assign BBM185=b[5]^b[12];
assign BBM186=b[0]^b[8];
assign BBM187=b[1]^b[9];
assign BBM188=b[3]^b[5];
assign BBM189=b[4]^b[7];
assign BBM190=b[4]^b[10];
assign BBM191=b[1]^b[8];
assign BBM192=b[6]^b[7];
assign BBM193=b[5]^b[9];
assign BBM194=b[8]^b[11];
assign BBM195=b[4]^b[9];
assign BBM196=b[3]^b[8];
assign BBM197=b[5]^b[11];
assign BBM198=b[10]^b[11];
assign BBM199=b[1]^b[11];
assign BBM200=b[1]^b[10];
assign BBM201=b[2]^b[5];
assign BBM202=b[8]^b[9];
assign BBM203=b[2]^b[3];
assign BBM204=b[2]^b[6];
assign BBM205=b[0]^b[10];
assign BBM206=b[4]^b[5];
assign BBM207=b[11]^b[12];
assign BBM208=b[2]^b[10];
assign BBM209=b[9]^b[11];
assign BBM210=b[0]^b[1];
assign BBM211=b[7]^b[8];
assign BBM212=b[4]^b[10];
assign BBM213=b[4]^b[6];
assign BBM214=b[0]^b[8];
assign BBM215=b[8]^b[10];
assign BBM216=b[1]^b[12];
assign BBM217=b[7]^b[9];
assign BBM218=b[7]^b[11];
assign BBM219=b[8]^b[11];
assign BBM220=b[7]^b[10];
assign BBM221=b[5]^b[6];
assign BBM222=b[1]^b[11];
assign BBM223=b[6]^b[7];
assign BBM224=b[1]^b[9];
assign BBM225=b[1]^b[12];
assign BBM226=b[0]^b[10];
assign BBM227=b[2]^b[5];
assign BBM228=b[4]^b[6];
assign BBM229=b[2]^b[3];
assign BBM230=b[3]^b[8];
assign BBM231=b[5];


assign P[1]=BBM161;
assign P[2]=BBM162;
assign P[3]=BBM129;
assign P[4]=BBM96;
assign P[5]=BBM97;
assign P[6]=BBM130^b[11];
assign P[7]=BBM98;
assign P[8]=BBM131^b[0];
assign P[9]=BBM163^b[11];
assign P[10]=BBM164^b[11];
assign P[11]=BBM165;
assign P[13]=BBM97;
assign P[14]=BBM132^b[8];
assign P[15]=BBM99;
assign P[16]=BBM65^b[6];
assign P[17]=BBM66;
assign P[18]=BBM100;
assign P[19]=BBM101^b[3];
assign P[20]=BBM67^b[9];
assign P[21]=BBM68^b[1];
assign P[22]=BBM102^b[3];
assign P[23]=BBM69;
assign P[24]=BBM103;
assign P[25]=BBM96;
assign P[26]=BBM100;
assign P[27]=BBM70^BBM166;
assign P[28]=BBM71^BBM167;
assign P[29]=BBM22^b[0];
assign P[30]=BBM10;
assign P[31]=BBM23;
assign P[32]=BBM24;
assign P[33]=BBM25;
assign P[34]=BBM71^b[12];
assign P[35]=BBM104^b[12];
assign P[36]=BBM133^b[4];
assign P[37]=BBM105;
assign P[38]=BBM66;
assign P[39]=BBM23;
assign P[40]=BBM11;
assign P[41]=BBM26^b[0];
assign P[42]=BBM68^b[3];
assign P[43]=BBM1;
assign P[44]=BBM2;
assign P[45]=BBM3^BBM168;
assign P[46]=BBM4^b[2];
assign P[47]=BBM5^b[3];
assign P[48]=BBM12^b[6];
assign P[49]=BBM13;
assign P[50]=BBM47^b[7];
assign P[51]=BBM10;
assign P[52]=BBM2;
assign P[53]=BBM106;
assign P[54]=BBM72;
assign P[55]=BBM48^b[11];
assign P[56]=BBM27;
assign P[57]=BBM14;
assign P[58]=BBM15^b[3];
assign P[59]=BBM49^BBM169;
assign P[60]=BBM28^b[2];
assign P[61]=BBM28^BBM167;
assign P[62]=BBM16^b[7];
assign P[63]=BBM3^b[7];
assign P[64]=BBM1;
assign P[65]=BBM14;
assign P[66]=BBM133;
assign P[67]=BBM134;
assign P[68]=BBM29^b[10];
assign P[69]=BBM50;
assign P[70]=BBM73;
assign P[71]=BBM107^b[3];
assign P[72]=BBM135^b[4];
assign P[73]=BBM108;
assign P[74]=BBM109^b[11];
assign P[75]=BBM51;
assign P[76]=BBM70^b[2];
assign P[77]=BBM27;
assign P[78]=BBM73;
assign P[79]=BBM74^b[8];
assign P[80]=BBM75;
assign P[81]=BBM30^BBM162;
assign P[82]=BBM31;
assign P[83]=BBM52;
assign P[84]=BBM106^BBM170;
assign P[85]=BBM76^b[8];
assign P[86]=BBM77^b[8];
assign P[87]=BBM97^b[3];
assign P[88]=BBM78^b[7];
assign P[89]=BBM79^BBM171;
assign P[90]=BBM50;
assign P[91]=BBM52;
assign P[92]=BBM32^b[10];
assign P[93]=BBM17;
assign P[94]=BBM76^b[3];
assign P[95]=BBM80;
assign P[96]=BBM81;
assign P[97]=BBM102^b[10];
assign P[98]=BBM53;
assign P[99]=BBM82^b[4];
assign P[100]=BBM136^BBM172;
assign P[101]=BBM83^b[3];
assign P[102]=BBM67^BBM166;
assign P[103]=BBM31;
assign P[104]=BBM81;
assign P[105]=BBM132^BBM137;
assign P[106]=BBM84^BBM173;
assign P[107]=BBM47^b[9];
assign P[108]=BBM33;
assign P[109]=BBM54;
assign P[110]=BBM111^b[9];
assign P[111]=BBM112^b[10];
assign P[112]=BBM85^b[9];
assign P[113]=BBM55^b[12];
assign P[114]=BBM86^b[11];
assign P[115]=BBM111^b[12];
assign P[116]=BBM80;
assign P[117]=BBM54;
assign P[118]=BBM138^BBM174;
assign P[119]=BBM113;
assign P[120]=BBM6;
assign P[121]=BBM175;
assign P[122]=BBM139;
assign P[123]=BBM140^b[6];
assign P[124]=BBM109^b[2];
assign P[125]=BBM111^b[1];
assign P[126]=BBM112^b[2];
assign P[127]=BBM115^b[3];
assign P[128]=BBM85^b[6];
assign P[129]=BBM33;
assign P[130]=BBM139;
assign P[131]=BBM176^b[1];
assign P[132]=BBM141;
assign P[133]=BBM116^b[4];
assign P[134]=BBM142;
assign P[135]=BBM130;
assign P[136]=BBM143;
assign P[137]=BBM131;
assign P[138]=BBM144;
assign P[139]=BBM117;
assign P[140]=BBM145;
assign P[141]=BBM177;
assign P[142]=BBM175;
assign P[143]=BBM130;
assign P[144]=BBM147^b[9];
assign P[145]=BBM118;
assign P[146]=BBM65^BBM178;
assign P[147]=BBM87;
assign P[148]=BBM88;
assign P[149]=BBM119^b[9];
assign P[150]=BBM120^b[1];
assign P[151]=BBM148^b[3];
assign P[152]=BBM121;
assign P[153]=BBM149;
assign P[154]=BBM150;
assign P[155]=BBM142;
assign P[156]=BBM88;
assign P[157]=BBM34^b[11];
assign P[158]=BBM30^b[10];
assign P[159]=BBM35^b[4];
assign P[160]=BBM18;
assign P[161]=BBM7;
assign P[162]=BBM22^BBM179;
assign P[163]=BBM19;
assign P[164]=BBM36;
assign P[165]=BBM89^b[9];
assign P[166]=BBM56;
assign P[167]=BBM90^b[6];
assign P[168]=BBM87;
assign P[169]=BBM7;
assign P[170]=BBM37^b[8];
assign P[171]=BBM57^b[5];
assign P[172]=BBM151^b[7];
assign P[173]=BBM8;
assign P[174]=BBM9;
assign P[175]=BBM38^BBM180;
assign P[176]=BBM12^BBM170;
assign P[177]=BBM15^BBM181;
assign P[178]=BBM6^b[10];
assign P[179]=BBM26^BBM182;
assign P[180]=BBM32^BBM183;
assign P[181]=BBM18;
assign P[182]=BBM9;
assign P[183]=BBM91^b[4];
assign P[184]=BBM122^b[1];
assign P[185]=BBM99^b[1];
assign P[186]=BBM20;
assign P[187]=BBM21;
assign P[188]=BBM35^b[9];
assign P[189]=BBM27^b[6]^b[12];
assign P[190]=BBM39^b[7];
assign P[191]=BBM29^b[6];
assign P[192]=BBM49^BBM184;
assign P[193]=BBM58^BBM163;
assign P[194]=BBM8;
assign P[195]=BBM21;
assign P[196]=BBM40^b[3];
assign P[197]=BBM89^BBM185;
assign P[198]=BBM16^b[11];
assign P[199]=BBM41^b[6];
assign P[200]=BBM13^b[0];
assign P[201]=BBM17^b[7];
assign P[202]=BBM19^b[1];
assign P[203]=BBM36^b[2];
assign P[204]=BBM38^b[6];
assign P[205]=BBM40^b[1];
assign P[206]=BBM42^b[6];
assign P[207]=BBM20;
assign P[0]=b[5];
assign P[12]=b[4];


assign P1[12:0]=P[12:0];
assign P2[12:0]=P[25:13];
assign P3[12:0]=P[38:26];
assign P4[12:0]=P[51:39];
assign P5[12:0]=P[64:52];
assign P6[12:0]=P[77:65];
assign P7[12:0]=P[90:78];
assign P8[12:0]=P[103:91];
assign P9[12:0]=P[116:104];
assign P10[12:0]=P[129:117];
assign P11[12:0]=P[142:130];
assign P12[12:0]=P[155:143];
assign P13[12:0]=P[168:156];
assign P14[12:0]=P[181:169];
assign P15[12:0]=P[194:182];
assign P16[12:0]=P[207:195];









endmodule
