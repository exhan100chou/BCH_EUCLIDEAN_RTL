
module degree_computation_3_DW01_dec_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n1, n2, n3, n4, n5;

  XOR2X1 U1 ( .A(A[4]), .B(n1), .Y(SUM[4]) );
  NOR2X1 U2 ( .A(A[3]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[3]), .B(n2), .Y(SUM[3]) );
  OAI21XL U4 ( .A0(n3), .A1(n4), .B0(n2), .Y(SUM[2]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[2]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[1]) );
  AOI21X1 U8 ( .A0(A[0]), .A1(A[1]), .B0(n3), .Y(n5) );
  NOR2X1 U9 ( .A(A[1]), .B(A[0]), .Y(n3) );
  INVX1 U10 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module degree_computation_3_DW01_dec_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n1, n2, n3, n4, n5;

  XOR2X1 U1 ( .A(A[4]), .B(n1), .Y(SUM[4]) );
  NOR2X1 U2 ( .A(A[3]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[3]), .B(n2), .Y(SUM[3]) );
  OAI21XL U4 ( .A0(n3), .A1(n4), .B0(n2), .Y(SUM[2]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[2]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[1]) );
  AOI21X1 U8 ( .A0(A[0]), .A1(A[1]), .B0(n3), .Y(n5) );
  NOR2X1 U9 ( .A(A[1]), .B(A[0]), .Y(n3) );
  INVX1 U10 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module degree_computation_2_DW01_dec_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n1, n2, n3, n4, n5;

  XOR2X1 U1 ( .A(A[4]), .B(n1), .Y(SUM[4]) );
  NOR2X1 U2 ( .A(A[3]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[3]), .B(n2), .Y(SUM[3]) );
  OAI21XL U4 ( .A0(n3), .A1(n4), .B0(n2), .Y(SUM[2]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[2]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[1]) );
  AOI21X1 U8 ( .A0(A[0]), .A1(A[1]), .B0(n3), .Y(n5) );
  NOR2X1 U9 ( .A(A[1]), .B(A[0]), .Y(n3) );
  INVX1 U10 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module degree_computation_2_DW01_dec_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n1, n2, n3, n4, n5;

  XOR2X1 U1 ( .A(A[4]), .B(n1), .Y(SUM[4]) );
  NOR2X1 U2 ( .A(A[3]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[3]), .B(n2), .Y(SUM[3]) );
  OAI21XL U4 ( .A0(n3), .A1(n4), .B0(n2), .Y(SUM[2]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[2]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[1]) );
  AOI21X1 U8 ( .A0(A[0]), .A1(A[1]), .B0(n3), .Y(n5) );
  NOR2X1 U9 ( .A(A[1]), .B(A[0]), .Y(n3) );
  INVX1 U10 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module degree_computation_1_DW01_dec_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n1, n2, n3, n4, n5;

  XOR2X1 U1 ( .A(A[4]), .B(n1), .Y(SUM[4]) );
  NOR2X1 U2 ( .A(A[3]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[3]), .B(n2), .Y(SUM[3]) );
  OAI21XL U4 ( .A0(n3), .A1(n4), .B0(n2), .Y(SUM[2]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[2]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[1]) );
  AOI21X1 U8 ( .A0(A[0]), .A1(A[1]), .B0(n3), .Y(n5) );
  NOR2X1 U9 ( .A(A[1]), .B(A[0]), .Y(n3) );
  INVX1 U10 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module degree_computation_1_DW01_dec_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n1, n2, n3, n4, n5;

  XOR2X1 U1 ( .A(A[4]), .B(n1), .Y(SUM[4]) );
  NOR2X1 U2 ( .A(A[3]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[3]), .B(n2), .Y(SUM[3]) );
  OAI21XL U4 ( .A0(n3), .A1(n4), .B0(n2), .Y(SUM[2]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[2]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[1]) );
  AOI21X1 U8 ( .A0(A[0]), .A1(A[1]), .B0(n3), .Y(n5) );
  NOR2X1 U9 ( .A(A[1]), .B(A[0]), .Y(n3) );
  INVX1 U10 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module degree_computation_0_DW01_dec_1 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n1, n2, n3, n4, n5;

  XOR2X1 U1 ( .A(A[4]), .B(n1), .Y(SUM[4]) );
  NOR2X1 U2 ( .A(A[3]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[3]), .B(n2), .Y(SUM[3]) );
  OAI21XL U4 ( .A0(n3), .A1(n4), .B0(n2), .Y(SUM[2]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[2]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[1]) );
  AOI21X1 U8 ( .A0(A[0]), .A1(A[1]), .B0(n3), .Y(n5) );
  NOR2X1 U9 ( .A(A[1]), .B(A[0]), .Y(n3) );
  INVX1 U10 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module degree_computation_0_DW01_dec_0 ( A, SUM );
  input [4:0] A;
  output [4:0] SUM;
  wire   n1, n2, n3, n4, n5;

  XOR2X1 U1 ( .A(A[4]), .B(n1), .Y(SUM[4]) );
  NOR2X1 U2 ( .A(A[3]), .B(n2), .Y(n1) );
  XNOR2X1 U3 ( .A(A[3]), .B(n2), .Y(SUM[3]) );
  OAI21XL U4 ( .A0(n3), .A1(n4), .B0(n2), .Y(SUM[2]) );
  NAND2X1 U5 ( .A(n3), .B(n4), .Y(n2) );
  INVX1 U6 ( .A(A[2]), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(SUM[1]) );
  AOI21X1 U8 ( .A0(A[0]), .A1(A[1]), .B0(n3), .Y(n5) );
  NOR2X1 U9 ( .A(A[1]), .B(A[0]), .Y(n3) );
  INVX1 U10 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module euclidean_4cells_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;
  wire   \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] ;

  ADDHXL U1_1_8 ( .A(A[8]), .B(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  XOR2X1 U1 ( .A(\carry[9] ), .B(A[9]), .Y(SUM[9]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module correct_module_4cells_p16_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;
  wire   \carry[9] , \carry[8] , \carry[7] , \carry[6] , \carry[5] ,
         \carry[4] , \carry[3] , \carry[2] ;

  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(\carry[2] ), .S(SUM[1]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  XOR2X1 U1 ( .A(\carry[9] ), .B(A[9]), .Y(SUM[9]) );
  INVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module mux_13_52 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n1), .Y(n4) );
  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(sel), .Y(n3) );
  INVX1 U5 ( .A(n8), .Y(out[12]) );
  AOI22X1 U6 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n3), .Y(n8) );
  INVX1 U7 ( .A(n6), .Y(out[10]) );
  AOI22X1 U8 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n3), .Y(n6) );
  INVX1 U9 ( .A(n18), .Y(out[9]) );
  AOI22X1 U10 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  INVX1 U11 ( .A(n17), .Y(out[8]) );
  AOI22X1 U12 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n4), .Y(n17) );
  INVX1 U13 ( .A(n15), .Y(out[7]) );
  AOI22X1 U14 ( .A0(a[7]), .A1(n2), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U15 ( .A(n14), .Y(out[6]) );
  AOI22X1 U16 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n14) );
  INVX1 U17 ( .A(n13), .Y(out[5]) );
  AOI22X1 U18 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n4), .Y(n13) );
  INVX1 U19 ( .A(n12), .Y(out[4]) );
  AOI22X1 U20 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U21 ( .A(n11), .Y(out[3]) );
  AOI22X1 U22 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n3), .Y(n11) );
  INVX1 U23 ( .A(n10), .Y(out[2]) );
  AOI22X1 U24 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n4), .Y(n10) );
  INVX1 U25 ( .A(n9), .Y(out[1]) );
  AOI22X1 U26 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n4), .Y(n9) );
  INVX1 U27 ( .A(n5), .Y(out[0]) );
  AOI22X1 U28 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n4), .Y(n5) );
  INVX1 U29 ( .A(n7), .Y(out[11]) );
  AOI22X1 U30 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n7) );
endmodule


module mux_13_51 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  INVX1 U1 ( .A(sel), .Y(n3) );
  INVX1 U2 ( .A(n2), .Y(n1) );
  INVX1 U3 ( .A(sel), .Y(n2) );
  INVX1 U4 ( .A(n7), .Y(out[12]) );
  AOI22X1 U5 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n2), .Y(n7) );
  INVX1 U6 ( .A(n6), .Y(out[11]) );
  AOI22X1 U7 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n6) );
  INVX1 U8 ( .A(n5), .Y(out[10]) );
  AOI22X1 U9 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n5) );
  INVX1 U10 ( .A(n17), .Y(out[9]) );
  AOI22X1 U11 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  INVX1 U12 ( .A(n15), .Y(out[8]) );
  AOI22X1 U13 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n15) );
  INVX1 U14 ( .A(n14), .Y(out[7]) );
  AOI22X1 U15 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n3), .Y(n14) );
  INVX1 U16 ( .A(n13), .Y(out[6]) );
  AOI22X1 U17 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n3), .Y(n13) );
  INVX1 U18 ( .A(n12), .Y(out[5]) );
  AOI22X1 U19 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n3), .Y(n12) );
  INVX1 U20 ( .A(n11), .Y(out[4]) );
  AOI22X1 U21 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n2), .Y(n11) );
  INVX1 U22 ( .A(n10), .Y(out[3]) );
  AOI22X1 U23 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n3), .Y(n10) );
  INVX1 U24 ( .A(n9), .Y(out[2]) );
  AOI22X1 U25 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n9) );
  INVX1 U26 ( .A(n8), .Y(out[1]) );
  AOI22X1 U27 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n3), .Y(n8) );
  INVX1 U28 ( .A(n4), .Y(out[0]) );
  AOI22X1 U29 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n3), .Y(n4) );
endmodule


module mux_13_50 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n2), .Y(n4) );
  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(sel), .Y(n3) );
  INVX1 U5 ( .A(n6), .Y(out[10]) );
  AOI22X1 U6 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n6) );
  INVX1 U7 ( .A(n7), .Y(out[11]) );
  AOI22X1 U8 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n7) );
  INVX1 U9 ( .A(n8), .Y(out[12]) );
  AOI22X1 U10 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n3), .Y(n8) );
  INVX1 U11 ( .A(n18), .Y(out[9]) );
  AOI22X1 U12 ( .A0(n2), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n18) );
  INVX1 U13 ( .A(n17), .Y(out[8]) );
  AOI22X1 U14 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n4), .Y(n17) );
  INVX1 U15 ( .A(n15), .Y(out[7]) );
  AOI22X1 U16 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n4), .Y(n15) );
  INVX1 U17 ( .A(n14), .Y(out[6]) );
  AOI22X1 U18 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n3), .Y(n14) );
  INVX1 U19 ( .A(n13), .Y(out[5]) );
  AOI22X1 U20 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n4), .Y(n13) );
  INVX1 U21 ( .A(n12), .Y(out[4]) );
  AOI22X1 U22 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U23 ( .A(n11), .Y(out[3]) );
  AOI22X1 U24 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n3), .Y(n11) );
  INVX1 U25 ( .A(n10), .Y(out[2]) );
  AOI22X1 U26 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n3), .Y(n10) );
  INVX1 U27 ( .A(n9), .Y(out[1]) );
  AOI22X1 U28 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n3), .Y(n9) );
  INVX1 U29 ( .A(n5), .Y(out[0]) );
  AOI22X1 U30 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n4), .Y(n5) );
endmodule


module mux_13_49 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n4), .Y(n2) );
  INVX1 U2 ( .A(sel), .Y(n4) );
  INVX1 U3 ( .A(sel), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n1) );
  INVX1 U5 ( .A(n9), .Y(out[1]) );
  AOI22X1 U6 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n9) );
  INVX1 U7 ( .A(n5), .Y(out[0]) );
  AOI22X1 U8 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n5) );
  INVX1 U9 ( .A(n18), .Y(out[9]) );
  AOI22X1 U10 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n18) );
  INVX1 U11 ( .A(n8), .Y(out[12]) );
  AOI22X1 U12 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n3), .Y(n8) );
  INVX1 U13 ( .A(n7), .Y(out[11]) );
  AOI22X1 U14 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n4), .Y(n7) );
  INVX1 U15 ( .A(n6), .Y(out[10]) );
  AOI22X1 U16 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n4), .Y(n6) );
  INVX1 U17 ( .A(n17), .Y(out[8]) );
  AOI22X1 U18 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n4), .Y(n17) );
  INVX1 U19 ( .A(n15), .Y(out[7]) );
  AOI22X1 U20 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U21 ( .A(n14), .Y(out[6]) );
  AOI22X1 U22 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n14) );
  INVX1 U23 ( .A(n13), .Y(out[5]) );
  AOI22X1 U24 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n4), .Y(n13) );
  INVX1 U25 ( .A(n12), .Y(out[4]) );
  AOI22X1 U26 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U27 ( .A(n11), .Y(out[3]) );
  AOI22X1 U28 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n4), .Y(n11) );
  INVX1 U29 ( .A(n10), .Y(out[2]) );
  AOI22X1 U30 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n3), .Y(n10) );
endmodule


module mux_13_48 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n34, n35, n36, n37, n38;

  INVX1 U1 ( .A(n38), .Y(out[6]) );
  INVX1 U2 ( .A(a[6]), .Y(n1) );
  INVX1 U3 ( .A(a[12]), .Y(n2) );
  INVXL U4 ( .A(a[9]), .Y(n15) );
  INVX1 U5 ( .A(a[3]), .Y(n5) );
  INVX1 U6 ( .A(b[5]), .Y(n10) );
  INVX1 U7 ( .A(a[8]), .Y(n13) );
  INVX1 U8 ( .A(a[10]), .Y(n17) );
  AOI2BB2X1 U9 ( .B0(b[6]), .B1(n4), .A0N(n1), .A1N(n4), .Y(n38) );
  INVX1 U10 ( .A(n35), .Y(out[12]) );
  INVX1 U11 ( .A(n36), .Y(out[1]) );
  MXI2X1 U12 ( .A(n9), .B(n10), .S0(n4), .Y(out[5]) );
  AOI2BB2X1 U13 ( .B0(b[12]), .B1(n4), .A0N(n2), .A1N(n4), .Y(n35) );
  INVXL U14 ( .A(n37), .Y(out[2]) );
  INVXL U15 ( .A(a[4]), .Y(n7) );
  INVXL U16 ( .A(a[5]), .Y(n9) );
  INVXL U17 ( .A(a[7]), .Y(n11) );
  INVXL U18 ( .A(a[11]), .Y(n19) );
  INVX1 U19 ( .A(n4), .Y(n3) );
  INVX1 U20 ( .A(sel), .Y(n4) );
  INVX1 U21 ( .A(b[10]), .Y(n18) );
  INVX1 U22 ( .A(b[8]), .Y(n14) );
  INVX1 U23 ( .A(b[4]), .Y(n8) );
  INVX1 U24 ( .A(b[7]), .Y(n12) );
  INVX1 U25 ( .A(b[3]), .Y(n6) );
  INVX1 U26 ( .A(b[9]), .Y(n16) );
  INVX1 U27 ( .A(b[11]), .Y(n21) );
  MXI2X1 U28 ( .A(n6), .B(n5), .S0(n3), .Y(out[3]) );
  MXI2X1 U29 ( .A(n8), .B(n7), .S0(n3), .Y(out[4]) );
  MXI2X1 U30 ( .A(n14), .B(n13), .S0(n3), .Y(out[8]) );
  MXI2X1 U31 ( .A(n16), .B(n15), .S0(n3), .Y(out[9]) );
  MXI2X1 U32 ( .A(n18), .B(n17), .S0(n3), .Y(out[10]) );
  MXI2X1 U33 ( .A(n21), .B(n19), .S0(n3), .Y(out[11]) );
  MXI2X1 U34 ( .A(n12), .B(n11), .S0(n3), .Y(out[7]) );
  INVX1 U35 ( .A(n34), .Y(out[0]) );
  AOI22X1 U36 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n4), .Y(n34) );
  AOI22X1 U37 ( .A0(a[1]), .A1(n3), .B0(b[1]), .B1(n4), .Y(n36) );
  AOI22X1 U38 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n4), .Y(n37) );
endmodule


module mux_13_47 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  AOI22XL U1 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n4), .Y(n5) );
  AOI22XL U2 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n4), .Y(n9) );
  AOI22XL U3 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n1), .Y(n11) );
  AOI22XL U4 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  AOI22XL U5 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n4), .Y(n13) );
  AOI22XL U6 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n4), .Y(n14) );
  AOI22XL U7 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n4), .Y(n6) );
  AOI22XL U8 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n4), .Y(n7) );
  AOI22XL U9 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n1), .Y(n8) );
  AOI22XL U10 ( .A0(a[8]), .A1(n3), .B0(b[8]), .B1(n4), .Y(n17) );
  AOI22XL U11 ( .A0(a[7]), .A1(n3), .B0(b[7]), .B1(n1), .Y(n15) );
  AOI22XL U12 ( .A0(n3), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  INVX1 U14 ( .A(n4), .Y(n3) );
  INVX1 U15 ( .A(sel), .Y(n4) );
  INVX1 U16 ( .A(sel), .Y(n1) );
  INVX1 U17 ( .A(n5), .Y(out[0]) );
  INVX1 U18 ( .A(n9), .Y(out[1]) );
  INVX1 U19 ( .A(n10), .Y(out[2]) );
  AOI22X1 U20 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n1), .Y(n10) );
  INVX1 U21 ( .A(n11), .Y(out[3]) );
  INVX1 U22 ( .A(n12), .Y(out[4]) );
  INVX1 U23 ( .A(n13), .Y(out[5]) );
  INVX1 U24 ( .A(n14), .Y(out[6]) );
  INVX1 U25 ( .A(n15), .Y(out[7]) );
  INVX1 U26 ( .A(n17), .Y(out[8]) );
  INVX1 U27 ( .A(n18), .Y(out[9]) );
  INVX1 U28 ( .A(n6), .Y(out[10]) );
  INVX1 U29 ( .A(n7), .Y(out[11]) );
  INVX1 U30 ( .A(n8), .Y(out[12]) );
endmodule


module mux_13_46 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n34, n35, n36, n37, n38;

  CLKINVXL U1 ( .A(a[5]), .Y(n9) );
  CLKINVXL U2 ( .A(a[10]), .Y(n17) );
  INVX1 U3 ( .A(a[1]), .Y(n1) );
  AOI2BB2X1 U4 ( .B0(b[1]), .B1(n4), .A0N(n1), .A1N(n4), .Y(n36) );
  INVX1 U5 ( .A(n36), .Y(out[1]) );
  INVX1 U6 ( .A(a[12]), .Y(n2) );
  INVX1 U7 ( .A(a[9]), .Y(n15) );
  INVX1 U8 ( .A(a[3]), .Y(n5) );
  INVX1 U9 ( .A(a[8]), .Y(n13) );
  INVX1 U10 ( .A(a[11]), .Y(n19) );
  INVX1 U11 ( .A(n38), .Y(out[6]) );
  INVX1 U12 ( .A(n35), .Y(out[12]) );
  CLKINVX2 U13 ( .A(b[5]), .Y(n10) );
  AOI2BB2X1 U14 ( .B0(b[12]), .B1(n4), .A0N(n2), .A1N(n4), .Y(n35) );
  INVXL U15 ( .A(n37), .Y(out[2]) );
  INVX1 U16 ( .A(n4), .Y(n3) );
  INVX1 U17 ( .A(b[10]), .Y(n18) );
  INVX1 U18 ( .A(sel), .Y(n4) );
  INVX1 U19 ( .A(b[4]), .Y(n8) );
  INVX1 U20 ( .A(b[8]), .Y(n14) );
  INVX1 U21 ( .A(b[11]), .Y(n21) );
  INVX1 U22 ( .A(b[7]), .Y(n12) );
  INVX1 U23 ( .A(b[3]), .Y(n6) );
  INVX1 U24 ( .A(b[9]), .Y(n16) );
  MXI2X1 U25 ( .A(n6), .B(n5), .S0(n3), .Y(out[3]) );
  MXI2X1 U26 ( .A(n8), .B(n7), .S0(n3), .Y(out[4]) );
  MXI2X1 U27 ( .A(n12), .B(n11), .S0(n3), .Y(out[7]) );
  MXI2X1 U28 ( .A(n14), .B(n13), .S0(n3), .Y(out[8]) );
  MXI2X1 U29 ( .A(n16), .B(n15), .S0(n3), .Y(out[9]) );
  MXI2X1 U30 ( .A(n18), .B(n17), .S0(n3), .Y(out[10]) );
  MXI2X1 U31 ( .A(n10), .B(n9), .S0(n3), .Y(out[5]) );
  MXI2X1 U32 ( .A(n21), .B(n19), .S0(n3), .Y(out[11]) );
  AOI22X1 U33 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n4), .Y(n37) );
  INVX1 U34 ( .A(n34), .Y(out[0]) );
  AOI22X1 U35 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n4), .Y(n34) );
  AOI22X1 U36 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n4), .Y(n38) );
  INVX1 U37 ( .A(a[4]), .Y(n7) );
  INVX1 U38 ( .A(a[7]), .Y(n11) );
endmodule


module mux_13_45 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  AOI22XL U1 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n2), .Y(n5) );
  AOI22XL U2 ( .A0(a[1]), .A1(n3), .B0(b[1]), .B1(n2), .Y(n9) );
  AOI22XL U3 ( .A0(a[3]), .A1(n3), .B0(b[3]), .B1(n2), .Y(n11) );
  AOI22XL U4 ( .A0(a[4]), .A1(n3), .B0(b[4]), .B1(n4), .Y(n12) );
  AOI22XL U5 ( .A0(a[5]), .A1(n3), .B0(b[5]), .B1(n4), .Y(n13) );
  AOI22XL U6 ( .A0(a[6]), .A1(n3), .B0(b[6]), .B1(n4), .Y(n14) );
  AOI22XL U7 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n2), .Y(n15) );
  AOI22XL U8 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n4), .Y(n17) );
  AOI22XL U9 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  AOI22XL U10 ( .A0(a[10]), .A1(n3), .B0(b[10]), .B1(n4), .Y(n6) );
  AOI22XL U11 ( .A0(a[11]), .A1(n3), .B0(b[11]), .B1(n2), .Y(n7) );
  AOI22XL U12 ( .A0(a[12]), .A1(n3), .B0(b[12]), .B1(n4), .Y(n8) );
  INVX1 U13 ( .A(n2), .Y(n3) );
  INVX1 U14 ( .A(n1), .Y(n4) );
  INVX1 U15 ( .A(n2), .Y(n1) );
  INVX1 U16 ( .A(sel), .Y(n2) );
  INVX1 U17 ( .A(n5), .Y(out[0]) );
  INVX1 U18 ( .A(n9), .Y(out[1]) );
  INVX1 U19 ( .A(n10), .Y(out[2]) );
  AOI22X1 U20 ( .A0(a[2]), .A1(n3), .B0(b[2]), .B1(n2), .Y(n10) );
  INVX1 U21 ( .A(n11), .Y(out[3]) );
  INVX1 U22 ( .A(n12), .Y(out[4]) );
  INVX1 U23 ( .A(n13), .Y(out[5]) );
  INVX1 U24 ( .A(n14), .Y(out[6]) );
  INVX1 U25 ( .A(n15), .Y(out[7]) );
  INVX1 U26 ( .A(n17), .Y(out[8]) );
  INVX1 U27 ( .A(n18), .Y(out[9]) );
  INVX1 U28 ( .A(n6), .Y(out[10]) );
  INVX1 U29 ( .A(n7), .Y(out[11]) );
  INVX1 U30 ( .A(n8), .Y(out[12]) );
endmodule


module mux_13_44 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n1), .Y(n4) );
  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(sel), .Y(n3) );
  INVX1 U5 ( .A(n6), .Y(out[10]) );
  AOI22X1 U6 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n3), .Y(n6) );
  INVX1 U7 ( .A(n18), .Y(out[9]) );
  AOI22X1 U8 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  INVX1 U9 ( .A(n17), .Y(out[8]) );
  AOI22X1 U10 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n4), .Y(n17) );
  INVX1 U11 ( .A(n15), .Y(out[7]) );
  AOI22X1 U12 ( .A0(a[7]), .A1(n2), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U13 ( .A(n14), .Y(out[6]) );
  AOI22X1 U14 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n4), .Y(n14) );
  INVX1 U15 ( .A(n13), .Y(out[5]) );
  AOI22X1 U16 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n4), .Y(n13) );
  INVX1 U17 ( .A(n12), .Y(out[4]) );
  AOI22X1 U18 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U19 ( .A(n11), .Y(out[3]) );
  AOI22X1 U20 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n3), .Y(n11) );
  INVX1 U21 ( .A(n10), .Y(out[2]) );
  AOI22X1 U22 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n4), .Y(n10) );
  INVX1 U23 ( .A(n9), .Y(out[1]) );
  AOI22X1 U24 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n4), .Y(n9) );
  INVX1 U25 ( .A(n5), .Y(out[0]) );
  AOI22X1 U26 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n4), .Y(n5) );
  INVX1 U27 ( .A(n8), .Y(out[12]) );
  AOI22X1 U28 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n3), .Y(n8) );
  INVX1 U29 ( .A(n7), .Y(out[11]) );
  AOI22X1 U30 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n3), .Y(n7) );
endmodule


module mux_13_43 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  INVX1 U1 ( .A(n1), .Y(n3) );
  INVX1 U2 ( .A(n2), .Y(n1) );
  INVX1 U3 ( .A(sel), .Y(n2) );
  INVX1 U4 ( .A(n6), .Y(out[11]) );
  AOI22X1 U5 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n6) );
  INVX1 U6 ( .A(n5), .Y(out[10]) );
  AOI22X1 U7 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n5) );
  INVX1 U8 ( .A(n17), .Y(out[9]) );
  AOI22X1 U9 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  INVX1 U10 ( .A(n15), .Y(out[8]) );
  AOI22X1 U11 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n15) );
  INVX1 U12 ( .A(n14), .Y(out[7]) );
  AOI22X1 U13 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n3), .Y(n14) );
  INVX1 U14 ( .A(n13), .Y(out[6]) );
  AOI22X1 U15 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n3), .Y(n13) );
  INVX1 U16 ( .A(n12), .Y(out[5]) );
  AOI22X1 U17 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n12) );
  INVX1 U18 ( .A(n11), .Y(out[4]) );
  AOI22X1 U19 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n2), .Y(n11) );
  INVX1 U20 ( .A(n10), .Y(out[3]) );
  AOI22X1 U21 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n3), .Y(n10) );
  INVX1 U22 ( .A(n9), .Y(out[2]) );
  AOI22X1 U23 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n3), .Y(n9) );
  INVX1 U24 ( .A(n8), .Y(out[1]) );
  AOI22X1 U25 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n8) );
  INVX1 U26 ( .A(n4), .Y(out[0]) );
  AOI22X1 U27 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n3), .Y(n4) );
  INVX1 U28 ( .A(n7), .Y(out[12]) );
  AOI22X1 U29 ( .A0(a[12]), .A1(sel), .B0(b[12]), .B1(n3), .Y(n7) );
endmodule


module mux_13_42 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n2), .Y(n4) );
  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(sel), .Y(n3) );
  INVX1 U5 ( .A(n18), .Y(out[9]) );
  AOI22X1 U6 ( .A0(n2), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n18) );
  INVX1 U7 ( .A(n17), .Y(out[8]) );
  AOI22X1 U8 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n3), .Y(n17) );
  INVX1 U9 ( .A(n15), .Y(out[7]) );
  AOI22X1 U10 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U11 ( .A(n14), .Y(out[6]) );
  AOI22X1 U12 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n3), .Y(n14) );
  INVX1 U13 ( .A(n13), .Y(out[5]) );
  AOI22X1 U14 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n3), .Y(n13) );
  INVX1 U15 ( .A(n12), .Y(out[4]) );
  AOI22X1 U16 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n3), .Y(n12) );
  INVX1 U17 ( .A(n11), .Y(out[3]) );
  AOI22X1 U18 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n3), .Y(n11) );
  INVX1 U19 ( .A(n10), .Y(out[2]) );
  AOI22X1 U20 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n4), .Y(n10) );
  INVX1 U21 ( .A(n9), .Y(out[1]) );
  AOI22X1 U22 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n4), .Y(n9) );
  INVX1 U23 ( .A(n5), .Y(out[0]) );
  AOI22X1 U24 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n4), .Y(n5) );
  INVX1 U25 ( .A(n8), .Y(out[12]) );
  AOI22X1 U26 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n4), .Y(n8) );
  INVX1 U27 ( .A(n7), .Y(out[11]) );
  AOI22X1 U28 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n4), .Y(n7) );
  INVX1 U29 ( .A(n6), .Y(out[10]) );
  AOI22X1 U30 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n6) );
endmodule


module mux_13_41 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n4), .Y(n2) );
  INVX1 U2 ( .A(sel), .Y(n4) );
  INVX1 U3 ( .A(sel), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(n1) );
  INVX1 U5 ( .A(n9), .Y(out[1]) );
  AOI22X1 U6 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n9) );
  INVX1 U7 ( .A(n5), .Y(out[0]) );
  AOI22X1 U8 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n5) );
  INVX1 U9 ( .A(n18), .Y(out[9]) );
  AOI22X1 U10 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n18) );
  INVX1 U11 ( .A(n8), .Y(out[12]) );
  AOI22X1 U12 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n3), .Y(n8) );
  INVX1 U13 ( .A(n7), .Y(out[11]) );
  AOI22X1 U14 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n4), .Y(n7) );
  INVX1 U15 ( .A(n6), .Y(out[10]) );
  AOI22X1 U16 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n4), .Y(n6) );
  INVX1 U17 ( .A(n17), .Y(out[8]) );
  AOI22X1 U18 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n4), .Y(n17) );
  INVX1 U19 ( .A(n15), .Y(out[7]) );
  AOI22X1 U20 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U21 ( .A(n14), .Y(out[6]) );
  AOI22X1 U22 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n14) );
  INVX1 U23 ( .A(n13), .Y(out[5]) );
  AOI22X1 U24 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n4), .Y(n13) );
  INVX1 U25 ( .A(n12), .Y(out[4]) );
  AOI22X1 U26 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U27 ( .A(n11), .Y(out[3]) );
  AOI22X1 U28 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n4), .Y(n11) );
  INVX1 U29 ( .A(n10), .Y(out[2]) );
  AOI22X1 U30 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n3), .Y(n10) );
endmodule


module mux_13_40 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n22, n35, n36, n37, n38, n39;

  INVXL U1 ( .A(a[9]), .Y(n16) );
  INVX1 U2 ( .A(n4), .Y(n2) );
  INVX1 U3 ( .A(a[1]), .Y(n1) );
  AOI2BB2X1 U4 ( .B0(b[1]), .B1(n5), .A0N(n1), .A1N(n2), .Y(n37) );
  INVX1 U5 ( .A(a[12]), .Y(n3) );
  INVX1 U6 ( .A(a[3]), .Y(n6) );
  INVX1 U7 ( .A(a[8]), .Y(n14) );
  MXI2X1 U8 ( .A(n10), .B(n11), .S0(n5), .Y(out[5]) );
  INVX1 U9 ( .A(n36), .Y(out[12]) );
  CLKINVX2 U10 ( .A(b[5]), .Y(n11) );
  AOI2BB2X1 U11 ( .B0(b[12]), .B1(n5), .A0N(n3), .A1N(n5), .Y(n36) );
  INVX1 U12 ( .A(a[10]), .Y(n18) );
  INVXL U13 ( .A(n38), .Y(out[2]) );
  INVXL U14 ( .A(n37), .Y(out[1]) );
  INVXL U15 ( .A(n39), .Y(out[6]) );
  INVXL U16 ( .A(a[4]), .Y(n8) );
  INVXL U17 ( .A(a[5]), .Y(n10) );
  INVXL U18 ( .A(a[7]), .Y(n12) );
  INVXL U19 ( .A(a[11]), .Y(n21) );
  INVX1 U20 ( .A(b[10]), .Y(n19) );
  INVX1 U21 ( .A(n5), .Y(n4) );
  INVX1 U22 ( .A(b[8]), .Y(n15) );
  INVX1 U23 ( .A(b[4]), .Y(n9) );
  INVX1 U24 ( .A(b[7]), .Y(n13) );
  INVX1 U25 ( .A(b[3]), .Y(n7) );
  INVX1 U26 ( .A(b[9]), .Y(n17) );
  INVX1 U27 ( .A(b[11]), .Y(n22) );
  INVX1 U28 ( .A(sel), .Y(n5) );
  MXI2X1 U29 ( .A(n9), .B(n8), .S0(n4), .Y(out[4]) );
  MXI2X1 U30 ( .A(n13), .B(n12), .S0(n4), .Y(out[7]) );
  MXI2X1 U31 ( .A(n7), .B(n6), .S0(n4), .Y(out[3]) );
  MXI2X1 U32 ( .A(n15), .B(n14), .S0(n4), .Y(out[8]) );
  MXI2X1 U33 ( .A(n17), .B(n16), .S0(n4), .Y(out[9]) );
  MXI2X1 U34 ( .A(n19), .B(n18), .S0(n4), .Y(out[10]) );
  MXI2X1 U35 ( .A(n22), .B(n21), .S0(n4), .Y(out[11]) );
  AOI22X1 U36 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n38) );
  INVX1 U37 ( .A(n35), .Y(out[0]) );
  AOI22X1 U38 ( .A0(a[0]), .A1(n4), .B0(b[0]), .B1(n5), .Y(n35) );
  AOI22X1 U39 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n5), .Y(n39) );
endmodule


module mux_13_39 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n1), .Y(n4) );
  AOI22XL U2 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n8) );
  AOI22XL U3 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n1), .Y(n9) );
  AOI22XL U4 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n1), .Y(n10) );
  AOI22XL U5 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n3), .Y(n11) );
  AOI22XL U6 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n3), .Y(n12) );
  AOI22XL U7 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n13) );
  AOI22XL U8 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n3), .Y(n14) );
  AOI22XL U9 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  AOI22XL U10 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n1), .Y(n7) );
  AOI22XL U11 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n3), .Y(n15) );
  AOI22XL U12 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n1), .Y(n6) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  INVX1 U14 ( .A(sel), .Y(n3) );
  INVX1 U15 ( .A(n4), .Y(out[0]) );
  INVX1 U16 ( .A(n8), .Y(out[1]) );
  INVX1 U17 ( .A(n9), .Y(out[2]) );
  INVX1 U18 ( .A(n10), .Y(out[3]) );
  INVX1 U19 ( .A(n11), .Y(out[4]) );
  INVX1 U20 ( .A(n12), .Y(out[5]) );
  INVX1 U21 ( .A(n13), .Y(out[6]) );
  INVX1 U22 ( .A(n14), .Y(out[7]) );
  INVX1 U23 ( .A(n15), .Y(out[8]) );
  INVX1 U24 ( .A(n17), .Y(out[9]) );
  INVX1 U25 ( .A(n5), .Y(out[10]) );
  AOI22X1 U26 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n3), .Y(n5) );
  INVX1 U27 ( .A(n6), .Y(out[11]) );
  INVX1 U28 ( .A(n7), .Y(out[12]) );
  INVX1 U29 ( .A(sel), .Y(n1) );
endmodule


module mux_13_38 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n33, n34, n35, n36, n37;

  INVX1 U1 ( .A(n35), .Y(out[1]) );
  INVXL U2 ( .A(n36), .Y(out[2]) );
  INVX1 U3 ( .A(n34), .Y(out[12]) );
  INVX1 U4 ( .A(a[12]), .Y(n1) );
  INVX1 U5 ( .A(a[3]), .Y(n4) );
  INVX1 U6 ( .A(a[8]), .Y(n12) );
  INVX1 U7 ( .A(a[11]), .Y(n18) );
  MXI2X1 U8 ( .A(n8), .B(n9), .S0(n3), .Y(out[5]) );
  AOI2BB2X1 U9 ( .B0(b[12]), .B1(n3), .A0N(n1), .A1N(n3), .Y(n34) );
  CLKINVX2 U10 ( .A(b[5]), .Y(n9) );
  INVX1 U11 ( .A(a[10]), .Y(n16) );
  INVXL U12 ( .A(n37), .Y(out[6]) );
  INVXL U13 ( .A(a[5]), .Y(n8) );
  INVXL U14 ( .A(a[9]), .Y(n14) );
  INVX1 U15 ( .A(b[10]), .Y(n17) );
  INVX1 U16 ( .A(n3), .Y(n2) );
  INVX1 U17 ( .A(b[11]), .Y(n19) );
  INVX1 U18 ( .A(b[8]), .Y(n13) );
  INVX1 U19 ( .A(b[7]), .Y(n11) );
  INVX1 U20 ( .A(b[3]), .Y(n5) );
  INVX1 U21 ( .A(b[4]), .Y(n7) );
  INVX1 U22 ( .A(b[9]), .Y(n15) );
  INVX1 U23 ( .A(sel), .Y(n3) );
  MXI2X1 U24 ( .A(n5), .B(n4), .S0(n2), .Y(out[3]) );
  MXI2X1 U25 ( .A(n7), .B(n6), .S0(n2), .Y(out[4]) );
  MXI2X1 U26 ( .A(n11), .B(n10), .S0(n2), .Y(out[7]) );
  MXI2X1 U27 ( .A(n13), .B(n12), .S0(n2), .Y(out[8]) );
  MXI2X1 U28 ( .A(n15), .B(n14), .S0(n2), .Y(out[9]) );
  MXI2X1 U29 ( .A(n17), .B(n16), .S0(n2), .Y(out[10]) );
  MXI2X1 U30 ( .A(n19), .B(n18), .S0(n2), .Y(out[11]) );
  INVX1 U31 ( .A(n33), .Y(out[0]) );
  AOI22X1 U32 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n33) );
  AOI22X1 U33 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n35) );
  AOI22X1 U34 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n3), .Y(n37) );
  AOI22X1 U35 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n3), .Y(n36) );
  INVX1 U36 ( .A(a[4]), .Y(n6) );
  INVX1 U37 ( .A(a[7]), .Y(n10) );
endmodule


module mux_13_37 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  AOI22XL U1 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n2), .Y(n5) );
  AOI22XL U2 ( .A0(a[1]), .A1(n3), .B0(b[1]), .B1(n4), .Y(n9) );
  AOI22XL U3 ( .A0(a[3]), .A1(n3), .B0(b[3]), .B1(n2), .Y(n11) );
  AOI22XL U4 ( .A0(a[4]), .A1(n3), .B0(b[4]), .B1(n4), .Y(n12) );
  AOI22XL U5 ( .A0(a[5]), .A1(n3), .B0(b[5]), .B1(n4), .Y(n13) );
  AOI22XL U6 ( .A0(a[6]), .A1(n3), .B0(b[6]), .B1(n2), .Y(n14) );
  AOI22XL U7 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n2), .Y(n15) );
  AOI22XL U8 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n17) );
  AOI22XL U9 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  AOI22XL U10 ( .A0(a[10]), .A1(n3), .B0(b[10]), .B1(n4), .Y(n6) );
  AOI22XL U11 ( .A0(a[11]), .A1(n3), .B0(b[11]), .B1(n2), .Y(n7) );
  AOI22XL U12 ( .A0(a[12]), .A1(n3), .B0(b[12]), .B1(n4), .Y(n8) );
  INVX1 U13 ( .A(n2), .Y(n3) );
  INVX1 U14 ( .A(n1), .Y(n4) );
  INVX1 U15 ( .A(n2), .Y(n1) );
  INVX1 U16 ( .A(sel), .Y(n2) );
  INVX1 U17 ( .A(n5), .Y(out[0]) );
  INVX1 U18 ( .A(n9), .Y(out[1]) );
  INVX1 U19 ( .A(n10), .Y(out[2]) );
  AOI22X1 U20 ( .A0(a[2]), .A1(n3), .B0(b[2]), .B1(n2), .Y(n10) );
  INVX1 U21 ( .A(n11), .Y(out[3]) );
  INVX1 U22 ( .A(n12), .Y(out[4]) );
  INVX1 U23 ( .A(n13), .Y(out[5]) );
  INVX1 U24 ( .A(n14), .Y(out[6]) );
  INVX1 U25 ( .A(n15), .Y(out[7]) );
  INVX1 U26 ( .A(n17), .Y(out[8]) );
  INVX1 U27 ( .A(n18), .Y(out[9]) );
  INVX1 U28 ( .A(n6), .Y(out[10]) );
  INVX1 U29 ( .A(n7), .Y(out[11]) );
  INVX1 U30 ( .A(n8), .Y(out[12]) );
endmodule


module mux_13_36 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n1), .Y(n4) );
  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(sel), .Y(n3) );
  INVX1 U5 ( .A(n6), .Y(out[10]) );
  AOI22X1 U6 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n4), .Y(n6) );
  INVX1 U7 ( .A(n18), .Y(out[9]) );
  AOI22X1 U8 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  INVX1 U9 ( .A(n17), .Y(out[8]) );
  AOI22X1 U10 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n4), .Y(n17) );
  INVX1 U11 ( .A(n15), .Y(out[7]) );
  AOI22X1 U12 ( .A0(a[7]), .A1(n2), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U13 ( .A(n14), .Y(out[6]) );
  AOI22X1 U14 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n14) );
  INVX1 U15 ( .A(n13), .Y(out[5]) );
  AOI22X1 U16 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n4), .Y(n13) );
  INVX1 U17 ( .A(n12), .Y(out[4]) );
  AOI22X1 U18 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U19 ( .A(n11), .Y(out[3]) );
  AOI22X1 U20 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n4), .Y(n11) );
  INVX1 U21 ( .A(n9), .Y(out[1]) );
  AOI22X1 U22 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n9) );
  INVX1 U23 ( .A(n5), .Y(out[0]) );
  AOI22X1 U24 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n4), .Y(n5) );
  INVX1 U25 ( .A(n10), .Y(out[2]) );
  AOI22X1 U26 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n4), .Y(n10) );
  INVX1 U27 ( .A(n8), .Y(out[12]) );
  AOI22X1 U28 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n3), .Y(n8) );
  INVX1 U29 ( .A(n7), .Y(out[11]) );
  AOI22X1 U30 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n7) );
endmodule


module mux_13_35 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  INVX1 U1 ( .A(sel), .Y(n3) );
  INVX1 U2 ( .A(n2), .Y(n1) );
  INVX1 U3 ( .A(sel), .Y(n2) );
  INVX1 U4 ( .A(n6), .Y(out[11]) );
  AOI22X1 U5 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n6) );
  INVX1 U6 ( .A(n5), .Y(out[10]) );
  AOI22X1 U7 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n2), .Y(n5) );
  INVX1 U8 ( .A(n17), .Y(out[9]) );
  AOI22X1 U9 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  INVX1 U10 ( .A(n15), .Y(out[8]) );
  AOI22X1 U11 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n15) );
  INVX1 U12 ( .A(n14), .Y(out[7]) );
  AOI22X1 U13 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n3), .Y(n14) );
  INVX1 U14 ( .A(n13), .Y(out[6]) );
  AOI22X1 U15 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n3), .Y(n13) );
  INVX1 U16 ( .A(n12), .Y(out[5]) );
  AOI22X1 U17 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n12) );
  INVX1 U18 ( .A(n11), .Y(out[4]) );
  AOI22X1 U19 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n3), .Y(n11) );
  INVX1 U20 ( .A(n10), .Y(out[3]) );
  AOI22X1 U21 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n3), .Y(n10) );
  INVX1 U22 ( .A(n8), .Y(out[1]) );
  AOI22X1 U23 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n3), .Y(n8) );
  INVX1 U24 ( .A(n4), .Y(out[0]) );
  AOI22X1 U25 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n3), .Y(n4) );
  INVX1 U26 ( .A(n7), .Y(out[12]) );
  AOI22X1 U27 ( .A0(a[12]), .A1(sel), .B0(b[12]), .B1(n3), .Y(n7) );
  INVX1 U28 ( .A(n9), .Y(out[2]) );
  AOI22X1 U29 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n9) );
endmodule


module mux_13_34 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n4), .Y(n2) );
  INVX1 U2 ( .A(sel), .Y(n3) );
  INVX1 U3 ( .A(sel), .Y(n4) );
  INVX1 U4 ( .A(n3), .Y(n1) );
  INVX1 U5 ( .A(n8), .Y(out[12]) );
  AOI22X1 U6 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n4), .Y(n8) );
  INVX1 U7 ( .A(n6), .Y(out[10]) );
  AOI22X1 U8 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n3), .Y(n6) );
  INVX1 U9 ( .A(n7), .Y(out[11]) );
  AOI22X1 U10 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n3), .Y(n7) );
  INVX1 U11 ( .A(n18), .Y(out[9]) );
  AOI22X1 U12 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n18) );
  INVX1 U13 ( .A(n17), .Y(out[8]) );
  AOI22X1 U14 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n3), .Y(n17) );
  INVX1 U15 ( .A(n15), .Y(out[7]) );
  AOI22X1 U16 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n4), .Y(n15) );
  INVX1 U17 ( .A(n14), .Y(out[6]) );
  AOI22X1 U18 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n4), .Y(n14) );
  INVX1 U19 ( .A(n13), .Y(out[5]) );
  AOI22X1 U20 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n3), .Y(n13) );
  INVX1 U21 ( .A(n12), .Y(out[4]) );
  AOI22X1 U22 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U23 ( .A(n11), .Y(out[3]) );
  AOI22X1 U24 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n4), .Y(n11) );
  INVX1 U25 ( .A(n10), .Y(out[2]) );
  AOI22X1 U26 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n3), .Y(n10) );
  INVX1 U27 ( .A(n9), .Y(out[1]) );
  AOI22X1 U28 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n4), .Y(n9) );
  INVX1 U29 ( .A(n5), .Y(out[0]) );
  AOI22X1 U30 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n5) );
endmodule


module mux_13_33 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n1), .Y(n4) );
  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(sel), .Y(n3) );
  INVX1 U5 ( .A(n9), .Y(out[1]) );
  AOI22X1 U6 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n3), .Y(n9) );
  INVX1 U7 ( .A(n5), .Y(out[0]) );
  AOI22X1 U8 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n5) );
  INVX1 U9 ( .A(n18), .Y(out[9]) );
  AOI22X1 U10 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  INVX1 U11 ( .A(n8), .Y(out[12]) );
  AOI22X1 U12 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n4), .Y(n8) );
  INVX1 U13 ( .A(n7), .Y(out[11]) );
  AOI22X1 U14 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n4), .Y(n7) );
  INVX1 U15 ( .A(n6), .Y(out[10]) );
  AOI22X1 U16 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n4), .Y(n6) );
  INVX1 U17 ( .A(n17), .Y(out[8]) );
  AOI22X1 U18 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n4), .Y(n17) );
  INVX1 U19 ( .A(n15), .Y(out[7]) );
  AOI22X1 U20 ( .A0(a[7]), .A1(n2), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U21 ( .A(n14), .Y(out[6]) );
  AOI22X1 U22 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n3), .Y(n14) );
  INVX1 U23 ( .A(n13), .Y(out[5]) );
  AOI22X1 U24 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n3), .Y(n13) );
  INVX1 U25 ( .A(n12), .Y(out[4]) );
  AOI22X1 U26 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U27 ( .A(n11), .Y(out[3]) );
  AOI22X1 U28 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n3), .Y(n11) );
  INVX1 U29 ( .A(n10), .Y(out[2]) );
  AOI22X1 U30 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n4), .Y(n10) );
endmodule


module mux_13_32 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n21, n34, n35, n36, n37, n38;

  INVX1 U1 ( .A(n37), .Y(out[2]) );
  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(a[1]), .Y(n1) );
  AOI2BB2X1 U4 ( .B0(b[1]), .B1(n4), .A0N(n1), .A1N(n2), .Y(n36) );
  INVXL U5 ( .A(a[9]), .Y(n15) );
  INVX1 U6 ( .A(a[3]), .Y(n5) );
  INVX1 U7 ( .A(a[8]), .Y(n13) );
  INVX1 U8 ( .A(n35), .Y(out[12]) );
  INVX1 U9 ( .A(n36), .Y(out[1]) );
  INVX1 U10 ( .A(n38), .Y(out[6]) );
  AOI22X1 U11 ( .A0(b[12]), .A1(n4), .B0(a[12]), .B1(sel), .Y(n35) );
  INVXL U12 ( .A(a[10]), .Y(n17) );
  MXI2X1 U13 ( .A(n9), .B(n10), .S0(n4), .Y(out[5]) );
  CLKINVX2 U14 ( .A(b[5]), .Y(n10) );
  INVXL U15 ( .A(a[4]), .Y(n7) );
  INVXL U16 ( .A(a[5]), .Y(n9) );
  INVXL U17 ( .A(a[7]), .Y(n11) );
  INVXL U18 ( .A(a[11]), .Y(n19) );
  INVX1 U19 ( .A(b[10]), .Y(n18) );
  INVX1 U20 ( .A(n4), .Y(n3) );
  INVX1 U21 ( .A(b[8]), .Y(n14) );
  INVX1 U22 ( .A(b[4]), .Y(n8) );
  INVX1 U23 ( .A(b[7]), .Y(n12) );
  INVX1 U24 ( .A(b[3]), .Y(n6) );
  INVX1 U25 ( .A(b[9]), .Y(n16) );
  INVX1 U26 ( .A(b[11]), .Y(n21) );
  INVX1 U27 ( .A(sel), .Y(n4) );
  MXI2X1 U28 ( .A(n12), .B(n11), .S0(n3), .Y(out[7]) );
  MXI2X1 U29 ( .A(n6), .B(n5), .S0(n3), .Y(out[3]) );
  MXI2X1 U30 ( .A(n8), .B(n7), .S0(n3), .Y(out[4]) );
  MXI2X1 U31 ( .A(n14), .B(n13), .S0(n3), .Y(out[8]) );
  MXI2X1 U32 ( .A(n16), .B(n15), .S0(n3), .Y(out[9]) );
  MXI2X1 U33 ( .A(n18), .B(n17), .S0(n3), .Y(out[10]) );
  MXI2X1 U34 ( .A(n21), .B(n19), .S0(n3), .Y(out[11]) );
  INVX1 U35 ( .A(n34), .Y(out[0]) );
  AOI22X1 U36 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n4), .Y(n34) );
  AOI22X1 U37 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n4), .Y(n38) );
  AOI22X1 U38 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n4), .Y(n37) );
endmodule


module mux_13_31 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n3), .Y(n15) );
  AOI22XL U2 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n3), .Y(n6) );
  AOI22XL U3 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n1), .Y(n4) );
  AOI22XL U4 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n1), .Y(n8) );
  AOI22XL U5 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n1), .Y(n10) );
  AOI22XL U6 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n3), .Y(n11) );
  AOI22XL U7 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n3), .Y(n12) );
  AOI22XL U8 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n13) );
  AOI22XL U9 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n3), .Y(n14) );
  AOI22XL U10 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  AOI22XL U11 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n1), .Y(n5) );
  AOI22XL U12 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n1), .Y(n7) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  INVX1 U14 ( .A(sel), .Y(n3) );
  INVX1 U15 ( .A(n4), .Y(out[0]) );
  INVX1 U16 ( .A(n8), .Y(out[1]) );
  INVX1 U17 ( .A(n9), .Y(out[2]) );
  AOI22X1 U18 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n3), .Y(n9) );
  INVX1 U19 ( .A(n10), .Y(out[3]) );
  INVX1 U20 ( .A(n11), .Y(out[4]) );
  INVX1 U21 ( .A(n12), .Y(out[5]) );
  INVX1 U22 ( .A(n13), .Y(out[6]) );
  INVX1 U23 ( .A(n14), .Y(out[7]) );
  INVX1 U24 ( .A(n15), .Y(out[8]) );
  INVX1 U25 ( .A(n17), .Y(out[9]) );
  INVX1 U26 ( .A(n5), .Y(out[10]) );
  INVX1 U27 ( .A(n6), .Y(out[11]) );
  INVX1 U28 ( .A(n7), .Y(out[12]) );
  INVX1 U29 ( .A(sel), .Y(n1) );
endmodule


module mux_13_30 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n33, n34, n35, n36, n37;

  INVXL U1 ( .A(n34), .Y(out[12]) );
  INVX1 U2 ( .A(a[12]), .Y(n1) );
  INVX1 U3 ( .A(a[3]), .Y(n4) );
  INVX1 U4 ( .A(a[8]), .Y(n12) );
  INVX1 U5 ( .A(a[11]), .Y(n18) );
  INVX1 U6 ( .A(n35), .Y(out[1]) );
  MXI2X1 U7 ( .A(n8), .B(n9), .S0(n3), .Y(out[5]) );
  AOI2BB2X1 U8 ( .B0(b[12]), .B1(n3), .A0N(n1), .A1N(n3), .Y(n34) );
  CLKINVX2 U9 ( .A(b[5]), .Y(n9) );
  INVX1 U10 ( .A(a[10]), .Y(n16) );
  INVXL U11 ( .A(n36), .Y(out[2]) );
  INVXL U12 ( .A(n37), .Y(out[6]) );
  INVXL U13 ( .A(a[5]), .Y(n8) );
  INVXL U14 ( .A(a[9]), .Y(n14) );
  INVX1 U15 ( .A(b[10]), .Y(n17) );
  INVX1 U16 ( .A(n3), .Y(n2) );
  INVX1 U17 ( .A(b[11]), .Y(n19) );
  INVX1 U18 ( .A(b[8]), .Y(n13) );
  INVX1 U19 ( .A(b[7]), .Y(n11) );
  INVX1 U20 ( .A(b[3]), .Y(n5) );
  INVX1 U21 ( .A(b[4]), .Y(n7) );
  INVX1 U22 ( .A(b[9]), .Y(n15) );
  INVX1 U23 ( .A(sel), .Y(n3) );
  MXI2X1 U24 ( .A(n5), .B(n4), .S0(n2), .Y(out[3]) );
  MXI2X1 U25 ( .A(n7), .B(n6), .S0(n2), .Y(out[4]) );
  MXI2X1 U26 ( .A(n11), .B(n10), .S0(n2), .Y(out[7]) );
  MXI2X1 U27 ( .A(n13), .B(n12), .S0(n2), .Y(out[8]) );
  MXI2X1 U28 ( .A(n15), .B(n14), .S0(n2), .Y(out[9]) );
  MXI2X1 U29 ( .A(n17), .B(n16), .S0(n2), .Y(out[10]) );
  MXI2X1 U30 ( .A(n19), .B(n18), .S0(n2), .Y(out[11]) );
  AOI22X1 U31 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n3), .Y(n36) );
  INVX1 U32 ( .A(n33), .Y(out[0]) );
  AOI22X1 U33 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n33) );
  AOI22X1 U34 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n35) );
  AOI22X1 U35 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n3), .Y(n37) );
  INVX1 U36 ( .A(a[4]), .Y(n6) );
  INVX1 U37 ( .A(a[7]), .Y(n10) );
endmodule


module mux_13_29 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n4) );
  AOI22XL U2 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n3), .Y(n8) );
  AOI22XL U3 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n2), .Y(n10) );
  AOI22XL U4 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n3), .Y(n11) );
  AOI22XL U5 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n3), .Y(n12) );
  AOI22XL U6 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n2), .Y(n13) );
  AOI22XL U7 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n2), .Y(n14) );
  AOI22XL U8 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n15) );
  AOI22XL U9 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  AOI22XL U10 ( .A0(a[10]), .A1(sel), .B0(b[10]), .B1(n3), .Y(n5) );
  AOI22XL U11 ( .A0(a[11]), .A1(sel), .B0(b[11]), .B1(n2), .Y(n6) );
  AOI22XL U12 ( .A0(a[12]), .A1(sel), .B0(b[12]), .B1(n3), .Y(n7) );
  INVX1 U13 ( .A(n1), .Y(n3) );
  INVX1 U14 ( .A(n2), .Y(n1) );
  INVX1 U15 ( .A(sel), .Y(n2) );
  INVX1 U16 ( .A(n4), .Y(out[0]) );
  INVX1 U17 ( .A(n8), .Y(out[1]) );
  INVX1 U18 ( .A(n9), .Y(out[2]) );
  AOI22X1 U19 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n9) );
  INVX1 U20 ( .A(n10), .Y(out[3]) );
  INVX1 U21 ( .A(n11), .Y(out[4]) );
  INVX1 U22 ( .A(n12), .Y(out[5]) );
  INVX1 U23 ( .A(n13), .Y(out[6]) );
  INVX1 U24 ( .A(n14), .Y(out[7]) );
  INVX1 U25 ( .A(n15), .Y(out[8]) );
  INVX1 U26 ( .A(n17), .Y(out[9]) );
  INVX1 U27 ( .A(n5), .Y(out[10]) );
  INVX1 U28 ( .A(n6), .Y(out[11]) );
  INVX1 U29 ( .A(n7), .Y(out[12]) );
endmodule


module mux_13_28 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n1), .Y(n4) );
  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(sel), .Y(n3) );
  INVX1 U5 ( .A(n7), .Y(out[11]) );
  AOI22X1 U6 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n7) );
  INVX1 U7 ( .A(n6), .Y(out[10]) );
  AOI22X1 U8 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n4), .Y(n6) );
  INVX1 U9 ( .A(n18), .Y(out[9]) );
  AOI22X1 U10 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  INVX1 U11 ( .A(n17), .Y(out[8]) );
  AOI22X1 U12 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n4), .Y(n17) );
  INVX1 U13 ( .A(n15), .Y(out[7]) );
  AOI22X1 U14 ( .A0(a[7]), .A1(n2), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U15 ( .A(n14), .Y(out[6]) );
  AOI22X1 U16 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n14) );
  INVX1 U17 ( .A(n13), .Y(out[5]) );
  AOI22X1 U18 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n3), .Y(n13) );
  INVX1 U19 ( .A(n12), .Y(out[4]) );
  AOI22X1 U20 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U21 ( .A(n11), .Y(out[3]) );
  AOI22X1 U22 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n3), .Y(n11) );
  INVX1 U23 ( .A(n10), .Y(out[2]) );
  AOI22X1 U24 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n4), .Y(n10) );
  INVX1 U25 ( .A(n9), .Y(out[1]) );
  AOI22X1 U26 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n9) );
  INVX1 U27 ( .A(n5), .Y(out[0]) );
  AOI22X1 U28 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n4), .Y(n5) );
  INVX1 U29 ( .A(n8), .Y(out[12]) );
  AOI22X1 U30 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n4), .Y(n8) );
endmodule


module mux_13_27 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  INVX1 U1 ( .A(n1), .Y(n3) );
  INVX1 U2 ( .A(n2), .Y(n1) );
  INVX1 U3 ( .A(sel), .Y(n2) );
  INVX1 U4 ( .A(n6), .Y(out[11]) );
  AOI22X1 U5 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n6) );
  INVX1 U6 ( .A(n5), .Y(out[10]) );
  AOI22X1 U7 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n5) );
  INVX1 U8 ( .A(n17), .Y(out[9]) );
  AOI22X1 U9 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  INVX1 U10 ( .A(n15), .Y(out[8]) );
  AOI22X1 U11 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n15) );
  INVX1 U12 ( .A(n14), .Y(out[7]) );
  AOI22X1 U13 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n3), .Y(n14) );
  INVX1 U14 ( .A(n13), .Y(out[6]) );
  AOI22X1 U15 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n3), .Y(n13) );
  INVX1 U16 ( .A(n12), .Y(out[5]) );
  AOI22X1 U17 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n12) );
  INVX1 U18 ( .A(n11), .Y(out[4]) );
  AOI22X1 U19 ( .A0(a[4]), .A1(sel), .B0(b[4]), .B1(n3), .Y(n11) );
  INVX1 U20 ( .A(n10), .Y(out[3]) );
  AOI22X1 U21 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n3), .Y(n10) );
  INVX1 U22 ( .A(n9), .Y(out[2]) );
  AOI22X1 U23 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n9) );
  INVX1 U24 ( .A(n8), .Y(out[1]) );
  AOI22X1 U25 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n8) );
  INVX1 U26 ( .A(n4), .Y(out[0]) );
  AOI22X1 U27 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n3), .Y(n4) );
  INVX1 U28 ( .A(n7), .Y(out[12]) );
  AOI22X1 U29 ( .A0(a[12]), .A1(sel), .B0(b[12]), .B1(n3), .Y(n7) );
endmodule


module mux_13_26 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n4), .Y(n2) );
  INVX1 U2 ( .A(sel), .Y(n3) );
  INVX1 U3 ( .A(sel), .Y(n4) );
  INVX1 U4 ( .A(n3), .Y(n1) );
  INVX1 U5 ( .A(n18), .Y(out[9]) );
  AOI22X1 U6 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n18) );
  INVX1 U7 ( .A(n17), .Y(out[8]) );
  AOI22X1 U8 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n4), .Y(n17) );
  INVX1 U9 ( .A(n15), .Y(out[7]) );
  AOI22X1 U10 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U11 ( .A(n14), .Y(out[6]) );
  AOI22X1 U12 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n14) );
  INVX1 U13 ( .A(n13), .Y(out[5]) );
  AOI22X1 U14 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n4), .Y(n13) );
  INVX1 U15 ( .A(n12), .Y(out[4]) );
  AOI22X1 U16 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U17 ( .A(n11), .Y(out[3]) );
  AOI22X1 U18 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n4), .Y(n11) );
  INVX1 U19 ( .A(n10), .Y(out[2]) );
  AOI22X1 U20 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n3), .Y(n10) );
  INVX1 U21 ( .A(n9), .Y(out[1]) );
  AOI22X1 U22 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n9) );
  INVX1 U23 ( .A(n5), .Y(out[0]) );
  AOI22X1 U24 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n5) );
  INVX1 U25 ( .A(n8), .Y(out[12]) );
  AOI22X1 U26 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n3), .Y(n8) );
  INVX1 U27 ( .A(n7), .Y(out[11]) );
  AOI22X1 U28 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n4), .Y(n7) );
  INVX1 U29 ( .A(n6), .Y(out[10]) );
  AOI22X1 U30 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n4), .Y(n6) );
endmodule


module mux_13_25 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n1), .Y(n4) );
  INVX1 U2 ( .A(n3), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(n1) );
  INVX1 U4 ( .A(sel), .Y(n3) );
  INVX1 U5 ( .A(n9), .Y(out[1]) );
  AOI22X1 U6 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n4), .Y(n9) );
  INVX1 U7 ( .A(n5), .Y(out[0]) );
  AOI22X1 U8 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n4), .Y(n5) );
  INVX1 U9 ( .A(n18), .Y(out[9]) );
  AOI22X1 U10 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  INVX1 U11 ( .A(n8), .Y(out[12]) );
  AOI22X1 U12 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n4), .Y(n8) );
  INVX1 U13 ( .A(n7), .Y(out[11]) );
  AOI22X1 U14 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n4), .Y(n7) );
  INVX1 U15 ( .A(n6), .Y(out[10]) );
  AOI22X1 U16 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n4), .Y(n6) );
  INVX1 U17 ( .A(n17), .Y(out[8]) );
  AOI22X1 U18 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n4), .Y(n17) );
  INVX1 U19 ( .A(n15), .Y(out[7]) );
  AOI22X1 U20 ( .A0(a[7]), .A1(n2), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U21 ( .A(n14), .Y(out[6]) );
  AOI22X1 U22 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n4), .Y(n14) );
  INVX1 U23 ( .A(n13), .Y(out[5]) );
  AOI22X1 U24 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n4), .Y(n13) );
  INVX1 U25 ( .A(n12), .Y(out[4]) );
  AOI22X1 U26 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n3), .Y(n12) );
  INVX1 U27 ( .A(n10), .Y(out[2]) );
  AOI22X1 U28 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n3), .Y(n10) );
  INVX1 U29 ( .A(n11), .Y(out[3]) );
  AOI22X1 U30 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n3), .Y(n11) );
endmodule


module mux_13_24 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n12, n13, n14, n15, n16;

  INVXL U1 ( .A(n13), .Y(out[12]) );
  INVXL U2 ( .A(a[12]), .Y(n1) );
  MX2XL U3 ( .A(b[9]), .B(a[9]), .S0(n2), .Y(out[9]) );
  AOI2BB2X1 U4 ( .B0(b[12]), .B1(n3), .A0N(n1), .A1N(n3), .Y(n13) );
  INVXL U5 ( .A(n15), .Y(out[2]) );
  INVXL U6 ( .A(n16), .Y(out[6]) );
  INVXL U7 ( .A(n14), .Y(out[1]) );
  INVX1 U8 ( .A(n3), .Y(n2) );
  INVX1 U9 ( .A(sel), .Y(n3) );
  MX2X1 U10 ( .A(b[5]), .B(a[5]), .S0(n2), .Y(out[5]) );
  MX2X1 U11 ( .A(b[7]), .B(a[7]), .S0(n2), .Y(out[7]) );
  MX2X1 U12 ( .A(b[3]), .B(a[3]), .S0(n2), .Y(out[3]) );
  MX2X1 U13 ( .A(b[11]), .B(a[11]), .S0(n2), .Y(out[11]) );
  MX2X1 U14 ( .A(b[10]), .B(a[10]), .S0(n2), .Y(out[10]) );
  MX2X1 U15 ( .A(b[8]), .B(a[8]), .S0(n2), .Y(out[8]) );
  MX2X1 U16 ( .A(b[4]), .B(a[4]), .S0(n2), .Y(out[4]) );
  AOI22X1 U17 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n3), .Y(n16) );
  AOI22X1 U18 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n3), .Y(n15) );
  AOI22X1 U19 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n14) );
  INVX1 U20 ( .A(n12), .Y(out[0]) );
  AOI22X1 U21 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n12) );
endmodule


module mux_13_23 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  AOI22XL U1 ( .A0(n3), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  AOI22XL U2 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n1), .Y(n9) );
  AOI22XL U3 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n1), .Y(n5) );
  AOI22XL U4 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n1), .Y(n8) );
  AOI22XL U5 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n1), .Y(n7) );
  AOI22XL U6 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n4), .Y(n14) );
  AOI22XL U7 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n4), .Y(n13) );
  AOI22XL U8 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n4), .Y(n12) );
  AOI22XL U9 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n1), .Y(n11) );
  AOI22XL U10 ( .A0(a[8]), .A1(n3), .B0(b[8]), .B1(n4), .Y(n17) );
  AOI22XL U11 ( .A0(a[7]), .A1(n3), .B0(b[7]), .B1(n4), .Y(n15) );
  INVX1 U12 ( .A(n1), .Y(n2) );
  INVX1 U13 ( .A(n4), .Y(n3) );
  INVX1 U14 ( .A(sel), .Y(n4) );
  INVX1 U15 ( .A(n18), .Y(out[9]) );
  INVX1 U16 ( .A(n8), .Y(out[12]) );
  INVX1 U17 ( .A(n7), .Y(out[11]) );
  INVX1 U18 ( .A(n6), .Y(out[10]) );
  AOI22X1 U19 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n4), .Y(n6) );
  INVX1 U20 ( .A(n14), .Y(out[6]) );
  INVX1 U21 ( .A(n13), .Y(out[5]) );
  INVX1 U22 ( .A(n12), .Y(out[4]) );
  INVX1 U23 ( .A(n11), .Y(out[3]) );
  INVX1 U24 ( .A(n10), .Y(out[2]) );
  AOI22X1 U25 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n1), .Y(n10) );
  INVX1 U26 ( .A(n9), .Y(out[1]) );
  INVX1 U27 ( .A(n5), .Y(out[0]) );
  INVX1 U28 ( .A(n17), .Y(out[8]) );
  INVX1 U29 ( .A(n15), .Y(out[7]) );
  INVX1 U30 ( .A(sel), .Y(n1) );
endmodule


module mux_13_22 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n12, n13, n14, n15, n16;

  MX2X2 U1 ( .A(b[3]), .B(a[3]), .S0(n2), .Y(out[3]) );
  INVX1 U2 ( .A(a[12]), .Y(n1) );
  MX2X2 U3 ( .A(b[5]), .B(a[5]), .S0(n2), .Y(out[5]) );
  AOI2BB2X1 U4 ( .B0(b[12]), .B1(n3), .A0N(n1), .A1N(n3), .Y(n13) );
  MX2X1 U5 ( .A(b[8]), .B(a[8]), .S0(n2), .Y(out[8]) );
  MX2X1 U6 ( .A(b[4]), .B(a[4]), .S0(n2), .Y(out[4]) );
  MX2X1 U7 ( .A(b[7]), .B(a[7]), .S0(n2), .Y(out[7]) );
  MX2X1 U8 ( .A(b[10]), .B(a[10]), .S0(n2), .Y(out[10]) );
  MX2X1 U9 ( .A(b[11]), .B(a[11]), .S0(n2), .Y(out[11]) );
  MX2X1 U10 ( .A(b[9]), .B(a[9]), .S0(n2), .Y(out[9]) );
  INVX1 U11 ( .A(n3), .Y(n2) );
  INVX1 U12 ( .A(sel), .Y(n3) );
  INVX1 U13 ( .A(n13), .Y(out[12]) );
  INVX1 U14 ( .A(n16), .Y(out[6]) );
  AOI22X1 U15 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n3), .Y(n16) );
  INVX1 U16 ( .A(n15), .Y(out[2]) );
  AOI22X1 U17 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n3), .Y(n15) );
  INVX1 U18 ( .A(n14), .Y(out[1]) );
  AOI22X1 U19 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n3), .Y(n14) );
  INVX1 U20 ( .A(n12), .Y(out[0]) );
  AOI22X1 U21 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n12) );
endmodule


module mux_13_21 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n4) );
  AOI22XL U2 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n3), .Y(n7) );
  AOI22XL U3 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n6) );
  AOI22XL U4 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n5) );
  AOI22XL U5 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n3), .Y(n13) );
  AOI22XL U6 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n12) );
  AOI22XL U7 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n2), .Y(n11) );
  AOI22XL U8 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n8) );
  AOI22XL U9 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n2), .Y(n15) );
  AOI22XL U10 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n2), .Y(n14) );
  AOI22XL U11 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n17) );
  INVX1 U12 ( .A(n3), .Y(n1) );
  INVX1 U13 ( .A(sel), .Y(n3) );
  INVX1 U14 ( .A(sel), .Y(n2) );
  INVX1 U15 ( .A(n10), .Y(out[3]) );
  INVX1 U16 ( .A(n9), .Y(out[2]) );
  INVX1 U17 ( .A(n7), .Y(out[12]) );
  INVX1 U18 ( .A(n6), .Y(out[11]) );
  INVX1 U19 ( .A(n5), .Y(out[10]) );
  INVX1 U20 ( .A(n13), .Y(out[6]) );
  INVX1 U21 ( .A(n12), .Y(out[5]) );
  INVX1 U22 ( .A(n11), .Y(out[4]) );
  INVX1 U23 ( .A(n8), .Y(out[1]) );
  INVX1 U24 ( .A(n4), .Y(out[0]) );
  INVX1 U25 ( .A(n17), .Y(out[9]) );
  INVX1 U26 ( .A(n15), .Y(out[8]) );
  INVX1 U27 ( .A(n14), .Y(out[7]) );
  AOI22X1 U28 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n9) );
  AOI22XL U29 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n3), .Y(n10) );
endmodule


module mux_13_20 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  INVX1 U1 ( .A(sel), .Y(n1) );
  BUFX3 U2 ( .A(n1), .Y(n3) );
  INVX1 U3 ( .A(n7), .Y(out[12]) );
  AOI22X1 U4 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n3), .Y(n7) );
  INVX1 U5 ( .A(n6), .Y(out[11]) );
  AOI22X1 U6 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n3), .Y(n6) );
  INVX1 U7 ( .A(n5), .Y(out[10]) );
  AOI22X1 U8 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n3), .Y(n5) );
  INVX1 U9 ( .A(n17), .Y(out[9]) );
  AOI22X1 U10 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  INVX1 U11 ( .A(n15), .Y(out[8]) );
  AOI22X1 U12 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n3), .Y(n15) );
  INVX1 U13 ( .A(n14), .Y(out[7]) );
  AOI22X1 U14 ( .A0(a[7]), .A1(n2), .B0(b[7]), .B1(n3), .Y(n14) );
  INVX1 U15 ( .A(n13), .Y(out[6]) );
  AOI22X1 U16 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n13) );
  INVX1 U17 ( .A(n12), .Y(out[5]) );
  AOI22X1 U18 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n3), .Y(n12) );
  INVX1 U19 ( .A(n11), .Y(out[4]) );
  AOI22X1 U20 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n3), .Y(n11) );
  INVX1 U21 ( .A(n10), .Y(out[3]) );
  AOI22X1 U22 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n1), .Y(n10) );
  INVX1 U23 ( .A(n9), .Y(out[2]) );
  AOI22X1 U24 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n1), .Y(n9) );
  INVX1 U25 ( .A(n8), .Y(out[1]) );
  AOI22X1 U26 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n1), .Y(n8) );
  INVX1 U27 ( .A(n4), .Y(out[0]) );
  AOI22X1 U28 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n3), .Y(n4) );
  BUFX3 U29 ( .A(sel), .Y(n2) );
endmodule


module mux_13_19 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n2), .Y(n13) );
  AOI22XL U2 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n14) );
  AOI22XL U3 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n17) );
  AOI22XL U4 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n15), .Y(n3) );
  AOI22XL U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n2), .Y(n9) );
  AOI22XL U6 ( .A0(a[12]), .A1(sel), .B0(b[12]), .B1(n15), .Y(n6) );
  AOI22XL U7 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n2), .Y(n12) );
  AOI22XL U8 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n7) );
  AOI22XL U9 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n11) );
  AOI22XL U10 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n2), .Y(n5) );
  AOI22XL U11 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n2), .Y(n10) );
  AOI22XL U12 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n2), .Y(n4) );
  INVX1 U13 ( .A(n17), .Y(out[9]) );
  INVX1 U14 ( .A(n14), .Y(out[8]) );
  INVX1 U15 ( .A(n13), .Y(out[7]) );
  BUFX3 U16 ( .A(n15), .Y(n2) );
  INVX1 U17 ( .A(n1), .Y(n15) );
  BUFX3 U18 ( .A(sel), .Y(n1) );
  INVX1 U19 ( .A(n12), .Y(out[6]) );
  INVX1 U20 ( .A(n9), .Y(out[3]) );
  INVX1 U21 ( .A(n6), .Y(out[12]) );
  INVX1 U22 ( .A(n3), .Y(out[0]) );
  INVX1 U23 ( .A(n11), .Y(out[5]) );
  INVX1 U24 ( .A(n8), .Y(out[2]) );
  AOI22X1 U25 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n15), .Y(n8) );
  INVX1 U26 ( .A(n5), .Y(out[11]) );
  INVX1 U27 ( .A(n10), .Y(out[4]) );
  INVX1 U28 ( .A(n7), .Y(out[1]) );
  INVX1 U29 ( .A(n4), .Y(out[10]) );
endmodule


module mux_13_18 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n3), .Y(n8) );
  AOI22XL U2 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n2), .Y(n7) );
  AOI22XL U3 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n6) );
  AOI22XL U4 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n5) );
  AOI22XL U5 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n3), .Y(n13) );
  AOI22XL U6 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n3), .Y(n12) );
  AOI22XL U7 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n3), .Y(n11) );
  AOI22XL U8 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n3), .Y(n10) );
  AOI22XL U9 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n3), .Y(n4) );
  AOI22XL U10 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n17) );
  AOI22XL U11 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n2), .Y(n15) );
  AOI22XL U12 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n2), .Y(n14) );
  INVX1 U13 ( .A(n2), .Y(n1) );
  INVX1 U14 ( .A(sel), .Y(n2) );
  INVX1 U15 ( .A(sel), .Y(n3) );
  INVX1 U16 ( .A(n7), .Y(out[12]) );
  INVX1 U17 ( .A(n6), .Y(out[11]) );
  INVX1 U18 ( .A(n5), .Y(out[10]) );
  INVX1 U19 ( .A(n17), .Y(out[9]) );
  INVX1 U20 ( .A(n15), .Y(out[8]) );
  INVX1 U21 ( .A(n14), .Y(out[7]) );
  INVX1 U22 ( .A(n13), .Y(out[6]) );
  INVX1 U23 ( .A(n12), .Y(out[5]) );
  INVX1 U24 ( .A(n11), .Y(out[4]) );
  INVX1 U25 ( .A(n10), .Y(out[3]) );
  INVX1 U26 ( .A(n9), .Y(out[2]) );
  AOI22X1 U27 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n3), .Y(n9) );
  INVX1 U28 ( .A(n8), .Y(out[1]) );
  INVX1 U29 ( .A(n4), .Y(out[0]) );
endmodule


module mux_13_17 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  AOI22XL U1 ( .A0(a[12]), .A1(n3), .B0(b[12]), .B1(n4), .Y(n8) );
  AOI22XL U2 ( .A0(a[10]), .A1(n3), .B0(b[10]), .B1(n2), .Y(n6) );
  AOI22XL U3 ( .A0(a[6]), .A1(n3), .B0(b[6]), .B1(n2), .Y(n14) );
  AOI22XL U4 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n18) );
  AOI22XL U5 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n2), .Y(n17) );
  AOI22XL U6 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n2), .Y(n15) );
  INVX1 U7 ( .A(n2), .Y(n3) );
  INVX1 U8 ( .A(n1), .Y(n4) );
  INVX1 U9 ( .A(n2), .Y(n1) );
  INVX1 U10 ( .A(sel), .Y(n2) );
  INVX1 U11 ( .A(n6), .Y(out[10]) );
  INVX1 U12 ( .A(n7), .Y(out[11]) );
  INVX1 U13 ( .A(n8), .Y(out[12]) );
  INVX1 U14 ( .A(n18), .Y(out[9]) );
  INVX1 U15 ( .A(n17), .Y(out[8]) );
  INVX1 U16 ( .A(n15), .Y(out[7]) );
  INVX1 U17 ( .A(n14), .Y(out[6]) );
  INVX1 U18 ( .A(n13), .Y(out[5]) );
  AOI22X1 U19 ( .A0(a[5]), .A1(n3), .B0(b[5]), .B1(n4), .Y(n13) );
  INVX1 U20 ( .A(n12), .Y(out[4]) );
  AOI22X1 U21 ( .A0(a[4]), .A1(n3), .B0(b[4]), .B1(n2), .Y(n12) );
  INVX1 U22 ( .A(n11), .Y(out[3]) );
  AOI22X1 U23 ( .A0(a[3]), .A1(n3), .B0(b[3]), .B1(n4), .Y(n11) );
  INVX1 U24 ( .A(n10), .Y(out[2]) );
  AOI22X1 U25 ( .A0(a[2]), .A1(n3), .B0(b[2]), .B1(n4), .Y(n10) );
  INVX1 U26 ( .A(n9), .Y(out[1]) );
  AOI22X1 U27 ( .A0(a[1]), .A1(n3), .B0(b[1]), .B1(n4), .Y(n9) );
  INVX1 U28 ( .A(n5), .Y(out[0]) );
  AOI22X1 U29 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n2), .Y(n5) );
  AOI22X1 U30 ( .A0(a[11]), .A1(n3), .B0(b[11]), .B1(n4), .Y(n7) );
endmodule


module mux_13_16 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  AOI22XL U1 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n3), .Y(n8) );
  AOI22XL U2 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n7) );
  AOI22XL U3 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n4), .Y(n6) );
  AOI22XL U4 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n3), .Y(n14) );
  AOI22XL U5 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n3), .Y(n12) );
  AOI22XL U6 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n4), .Y(n9) );
  AOI22XL U7 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n3), .Y(n5) );
  AOI22XL U8 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n3), .Y(n17) );
  AOI22XL U9 ( .A0(a[7]), .A1(n2), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U10 ( .A(n4), .Y(n1) );
  INVX1 U11 ( .A(n3), .Y(n2) );
  INVX1 U12 ( .A(sel), .Y(n3) );
  INVX1 U13 ( .A(sel), .Y(n4) );
  INVX1 U14 ( .A(n8), .Y(out[12]) );
  INVX1 U15 ( .A(n7), .Y(out[11]) );
  INVX1 U16 ( .A(n6), .Y(out[10]) );
  INVX1 U17 ( .A(n18), .Y(out[9]) );
  AOI22X1 U18 ( .A0(n2), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n18) );
  INVX1 U19 ( .A(n17), .Y(out[8]) );
  INVX1 U20 ( .A(n15), .Y(out[7]) );
  INVX1 U21 ( .A(n14), .Y(out[6]) );
  INVX1 U22 ( .A(n13), .Y(out[5]) );
  AOI22X1 U23 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n3), .Y(n13) );
  INVX1 U24 ( .A(n12), .Y(out[4]) );
  INVX1 U25 ( .A(n11), .Y(out[3]) );
  AOI22X1 U26 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n4), .Y(n11) );
  INVX1 U27 ( .A(n10), .Y(out[2]) );
  AOI22X1 U28 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n4), .Y(n10) );
  INVX1 U29 ( .A(n9), .Y(out[1]) );
  INVX1 U30 ( .A(n5), .Y(out[0]) );
endmodule


module mux_13_15 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n3), .Y(n7) );
  AOI22XL U2 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n3), .Y(n6) );
  AOI22XL U3 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n3), .Y(n5) );
  AOI22XL U4 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n1), .Y(n17) );
  AOI22XL U5 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n3), .Y(n15) );
  AOI22XL U6 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n1), .Y(n14) );
  INVX1 U7 ( .A(n1), .Y(n2) );
  INVX1 U8 ( .A(sel), .Y(n3) );
  INVX1 U9 ( .A(sel), .Y(n1) );
  INVX1 U10 ( .A(n7), .Y(out[12]) );
  INVX1 U11 ( .A(n6), .Y(out[11]) );
  INVX1 U12 ( .A(n5), .Y(out[10]) );
  INVX1 U13 ( .A(n17), .Y(out[9]) );
  INVX1 U14 ( .A(n15), .Y(out[8]) );
  INVX1 U15 ( .A(n14), .Y(out[7]) );
  INVX1 U16 ( .A(n13), .Y(out[6]) );
  AOI22X1 U17 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n13) );
  INVX1 U18 ( .A(n12), .Y(out[5]) );
  AOI22X1 U19 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n3), .Y(n12) );
  INVX1 U20 ( .A(n11), .Y(out[4]) );
  AOI22X1 U21 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n3), .Y(n11) );
  INVX1 U22 ( .A(n10), .Y(out[3]) );
  AOI22X1 U23 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n3), .Y(n10) );
  INVX1 U24 ( .A(n9), .Y(out[2]) );
  AOI22X1 U25 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n3), .Y(n9) );
  INVX1 U26 ( .A(n8), .Y(out[1]) );
  AOI22X1 U27 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n1), .Y(n8) );
  INVX1 U28 ( .A(n4), .Y(out[0]) );
  AOI22X1 U29 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n4) );
endmodule


module mux_13_14 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n2), .Y(n13) );
  AOI22XL U2 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n14) );
  AOI22XL U3 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n17) );
  AOI22XL U4 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n15), .Y(n3) );
  AOI22XL U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n2), .Y(n9) );
  AOI22XL U6 ( .A0(a[12]), .A1(sel), .B0(b[12]), .B1(n15), .Y(n6) );
  AOI22XL U7 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n2), .Y(n12) );
  AOI22XL U8 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n7) );
  AOI22XL U9 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n11) );
  AOI22XL U10 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n2), .Y(n5) );
  AOI22XL U11 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n2), .Y(n10) );
  AOI22XL U12 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n2), .Y(n4) );
  INVX1 U13 ( .A(n17), .Y(out[9]) );
  INVX1 U14 ( .A(n14), .Y(out[8]) );
  INVX1 U15 ( .A(n13), .Y(out[7]) );
  BUFX3 U16 ( .A(n15), .Y(n2) );
  INVX1 U17 ( .A(n1), .Y(n15) );
  BUFX3 U18 ( .A(sel), .Y(n1) );
  INVX1 U19 ( .A(n12), .Y(out[6]) );
  INVX1 U20 ( .A(n9), .Y(out[3]) );
  INVX1 U21 ( .A(n6), .Y(out[12]) );
  INVX1 U22 ( .A(n3), .Y(out[0]) );
  INVX1 U23 ( .A(n11), .Y(out[5]) );
  INVX1 U24 ( .A(n8), .Y(out[2]) );
  AOI22X1 U25 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n15), .Y(n8) );
  INVX1 U26 ( .A(n5), .Y(out[11]) );
  INVX1 U27 ( .A(n10), .Y(out[4]) );
  INVX1 U28 ( .A(n7), .Y(out[1]) );
  INVX1 U29 ( .A(n4), .Y(out[10]) );
endmodule


module mux_13_13 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n8) );
  AOI22XL U2 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n3), .Y(n7) );
  AOI22XL U3 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n3), .Y(n6) );
  AOI22XL U4 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n3), .Y(n5) );
  AOI22XL U5 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n1), .Y(n13) );
  AOI22XL U6 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n1), .Y(n12) );
  AOI22XL U7 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n1), .Y(n11) );
  AOI22XL U8 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n3), .Y(n10) );
  AOI22XL U9 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n1), .Y(n4) );
  AOI22XL U10 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n1), .Y(n17) );
  AOI22XL U11 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n1), .Y(n15) );
  AOI22XL U12 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n3), .Y(n14) );
  INVX1 U13 ( .A(n1), .Y(n2) );
  INVX1 U14 ( .A(sel), .Y(n3) );
  INVX1 U15 ( .A(n7), .Y(out[12]) );
  INVX1 U16 ( .A(n6), .Y(out[11]) );
  INVX1 U17 ( .A(n5), .Y(out[10]) );
  INVX1 U18 ( .A(n17), .Y(out[9]) );
  INVX1 U19 ( .A(n15), .Y(out[8]) );
  INVX1 U20 ( .A(n14), .Y(out[7]) );
  INVX1 U21 ( .A(n13), .Y(out[6]) );
  INVX1 U22 ( .A(n12), .Y(out[5]) );
  INVX1 U23 ( .A(n11), .Y(out[4]) );
  INVX1 U24 ( .A(n10), .Y(out[3]) );
  INVX1 U25 ( .A(n9), .Y(out[2]) );
  AOI22X1 U26 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n3), .Y(n9) );
  INVX1 U27 ( .A(n8), .Y(out[1]) );
  INVX1 U28 ( .A(n4), .Y(out[0]) );
  INVX1 U29 ( .A(sel), .Y(n1) );
endmodule


module mux_13_12 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  AOI22XL U1 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n4), .Y(n7) );
  AOI22XL U2 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n6) );
  AOI22XL U3 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n3), .Y(n14) );
  AOI22XL U4 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n3), .Y(n13) );
  AOI22XL U5 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n3), .Y(n12) );
  AOI22XL U6 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n4), .Y(n11) );
  AOI22XL U7 ( .A0(n2), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n18) );
  AOI22XL U8 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n3), .Y(n17) );
  AOI22XL U9 ( .A0(a[7]), .A1(n2), .B0(b[7]), .B1(n3), .Y(n15) );
  INVX1 U10 ( .A(n4), .Y(n1) );
  INVX1 U11 ( .A(n3), .Y(n2) );
  INVX1 U12 ( .A(sel), .Y(n3) );
  INVX1 U13 ( .A(sel), .Y(n4) );
  INVX1 U14 ( .A(n9), .Y(out[1]) );
  AOI22X1 U15 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n4), .Y(n9) );
  INVX1 U16 ( .A(n8), .Y(out[12]) );
  INVX1 U17 ( .A(n7), .Y(out[11]) );
  INVX1 U18 ( .A(n6), .Y(out[10]) );
  INVX1 U19 ( .A(n18), .Y(out[9]) );
  INVX1 U20 ( .A(n17), .Y(out[8]) );
  INVX1 U21 ( .A(n15), .Y(out[7]) );
  INVX1 U22 ( .A(n14), .Y(out[6]) );
  INVX1 U23 ( .A(n13), .Y(out[5]) );
  INVX1 U24 ( .A(n12), .Y(out[4]) );
  INVX1 U25 ( .A(n11), .Y(out[3]) );
  INVX1 U26 ( .A(n10), .Y(out[2]) );
  AOI22X1 U27 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n3), .Y(n10) );
  INVX1 U28 ( .A(n5), .Y(out[0]) );
  AOI22X1 U29 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n4), .Y(n5) );
  AOI22XL U30 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n4), .Y(n8) );
endmodule


module mux_13_11 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  AOI22XL U1 ( .A0(a[12]), .A1(n3), .B0(b[12]), .B1(n4), .Y(n8) );
  AOI22XL U2 ( .A0(a[10]), .A1(n3), .B0(b[10]), .B1(n2), .Y(n6) );
  AOI22XL U3 ( .A0(a[6]), .A1(n3), .B0(b[6]), .B1(n4), .Y(n14) );
  AOI22XL U4 ( .A0(a[4]), .A1(n3), .B0(b[4]), .B1(n4), .Y(n12) );
  AOI22XL U5 ( .A0(a[1]), .A1(n3), .B0(b[1]), .B1(n4), .Y(n9) );
  AOI22XL U6 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n2), .Y(n5) );
  AOI22XL U7 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n2), .Y(n17) );
  AOI22XL U8 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n4), .Y(n15) );
  INVX1 U9 ( .A(n2), .Y(n3) );
  INVX1 U10 ( .A(n1), .Y(n4) );
  INVX1 U11 ( .A(n2), .Y(n1) );
  INVX1 U12 ( .A(sel), .Y(n2) );
  INVX1 U13 ( .A(n8), .Y(out[12]) );
  INVX1 U14 ( .A(n7), .Y(out[11]) );
  AOI22X1 U15 ( .A0(a[11]), .A1(n3), .B0(b[11]), .B1(n2), .Y(n7) );
  INVX1 U16 ( .A(n6), .Y(out[10]) );
  INVX1 U17 ( .A(n18), .Y(out[9]) );
  AOI22X1 U18 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n18) );
  INVX1 U19 ( .A(n17), .Y(out[8]) );
  INVX1 U20 ( .A(n15), .Y(out[7]) );
  INVX1 U21 ( .A(n14), .Y(out[6]) );
  INVX1 U22 ( .A(n13), .Y(out[5]) );
  AOI22X1 U23 ( .A0(a[5]), .A1(n3), .B0(b[5]), .B1(n4), .Y(n13) );
  INVX1 U24 ( .A(n12), .Y(out[4]) );
  INVX1 U25 ( .A(n11), .Y(out[3]) );
  AOI22X1 U26 ( .A0(a[3]), .A1(n3), .B0(b[3]), .B1(n2), .Y(n11) );
  INVX1 U27 ( .A(n10), .Y(out[2]) );
  AOI22X1 U28 ( .A0(a[2]), .A1(n3), .B0(b[2]), .B1(n2), .Y(n10) );
  INVX1 U29 ( .A(n9), .Y(out[1]) );
  INVX1 U30 ( .A(n5), .Y(out[0]) );
endmodule


module mux_13_10 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n15) );
  AOI22XL U2 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n2), .Y(n7) );
  AOI22XL U3 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n2), .Y(n5) );
  AOI22XL U4 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n17) );
  AOI22XL U5 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n2), .Y(n14) );
  INVX1 U6 ( .A(n1), .Y(n3) );
  INVX1 U7 ( .A(n2), .Y(n1) );
  INVX1 U8 ( .A(sel), .Y(n2) );
  INVX1 U9 ( .A(n5), .Y(out[10]) );
  INVX1 U10 ( .A(n6), .Y(out[11]) );
  INVX1 U11 ( .A(n7), .Y(out[12]) );
  INVX1 U12 ( .A(n17), .Y(out[9]) );
  INVX1 U13 ( .A(n15), .Y(out[8]) );
  INVX1 U14 ( .A(n14), .Y(out[7]) );
  INVX1 U15 ( .A(n13), .Y(out[6]) );
  AOI22X1 U16 ( .A0(a[6]), .A1(sel), .B0(b[6]), .B1(n3), .Y(n13) );
  INVX1 U17 ( .A(n12), .Y(out[5]) );
  AOI22X1 U18 ( .A0(a[5]), .A1(sel), .B0(b[5]), .B1(n2), .Y(n12) );
  INVX1 U19 ( .A(n11), .Y(out[4]) );
  AOI22X1 U20 ( .A0(a[4]), .A1(sel), .B0(b[4]), .B1(n2), .Y(n11) );
  INVX1 U21 ( .A(n10), .Y(out[3]) );
  AOI22X1 U22 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n3), .Y(n10) );
  INVX1 U23 ( .A(n9), .Y(out[2]) );
  AOI22X1 U24 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n3), .Y(n9) );
  INVX1 U25 ( .A(n8), .Y(out[1]) );
  AOI22X1 U26 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n2), .Y(n8) );
  INVX1 U27 ( .A(n4), .Y(out[0]) );
  AOI22X1 U28 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n3), .Y(n4) );
  AOI22X1 U29 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n6) );
endmodule


module mux_13_9 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n2), .Y(n13) );
  AOI22XL U2 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n14) );
  AOI22XL U3 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n17) );
  AOI22XL U4 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n15), .Y(n3) );
  AOI22XL U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n2), .Y(n9) );
  AOI22XL U6 ( .A0(a[12]), .A1(sel), .B0(b[12]), .B1(n15), .Y(n6) );
  AOI22XL U7 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n2), .Y(n12) );
  AOI22XL U8 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n7) );
  AOI22XL U9 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n11) );
  AOI22XL U10 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n2), .Y(n5) );
  AOI22XL U11 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n2), .Y(n10) );
  AOI22XL U12 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n2), .Y(n4) );
  INVX1 U13 ( .A(n17), .Y(out[9]) );
  INVX1 U14 ( .A(n14), .Y(out[8]) );
  INVX1 U15 ( .A(n13), .Y(out[7]) );
  BUFX3 U16 ( .A(n15), .Y(n2) );
  INVX1 U17 ( .A(n1), .Y(n15) );
  BUFX3 U18 ( .A(sel), .Y(n1) );
  INVX1 U19 ( .A(n12), .Y(out[6]) );
  INVX1 U20 ( .A(n9), .Y(out[3]) );
  INVX1 U21 ( .A(n6), .Y(out[12]) );
  INVX1 U22 ( .A(n3), .Y(out[0]) );
  INVX1 U23 ( .A(n11), .Y(out[5]) );
  INVX1 U24 ( .A(n8), .Y(out[2]) );
  AOI22X1 U25 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n15), .Y(n8) );
  INVX1 U26 ( .A(n5), .Y(out[11]) );
  INVX1 U27 ( .A(n10), .Y(out[4]) );
  INVX1 U28 ( .A(n7), .Y(out[1]) );
  INVX1 U29 ( .A(n4), .Y(out[10]) );
endmodule


module mux_13_8 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n3), .Y(n8) );
  AOI22XL U2 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n3), .Y(n7) );
  AOI22XL U3 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n6) );
  AOI22XL U4 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n5) );
  AOI22XL U5 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n3), .Y(n13) );
  AOI22XL U6 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n3), .Y(n12) );
  AOI22XL U7 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n3), .Y(n11) );
  AOI22XL U8 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n3), .Y(n10) );
  AOI22XL U9 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n4) );
  AOI22XL U10 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n17) );
  AOI22XL U11 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n2), .Y(n15) );
  AOI22XL U12 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n2), .Y(n14) );
  INVX1 U13 ( .A(n2), .Y(n1) );
  INVX1 U14 ( .A(sel), .Y(n2) );
  INVX1 U15 ( .A(sel), .Y(n3) );
  INVX1 U16 ( .A(n7), .Y(out[12]) );
  INVX1 U17 ( .A(n6), .Y(out[11]) );
  INVX1 U18 ( .A(n5), .Y(out[10]) );
  INVX1 U19 ( .A(n17), .Y(out[9]) );
  INVX1 U20 ( .A(n15), .Y(out[8]) );
  INVX1 U21 ( .A(n14), .Y(out[7]) );
  INVX1 U22 ( .A(n13), .Y(out[6]) );
  INVX1 U23 ( .A(n12), .Y(out[5]) );
  INVX1 U24 ( .A(n11), .Y(out[4]) );
  INVX1 U25 ( .A(n10), .Y(out[3]) );
  INVX1 U26 ( .A(n9), .Y(out[2]) );
  AOI22X1 U27 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n3), .Y(n9) );
  INVX1 U28 ( .A(n8), .Y(out[1]) );
  INVX1 U29 ( .A(n4), .Y(out[0]) );
endmodule


module mux_13_7 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  AOI22XL U1 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n4), .Y(n17) );
  AOI22XL U2 ( .A0(a[10]), .A1(n3), .B0(b[10]), .B1(n4), .Y(n6) );
  AOI22XL U3 ( .A0(a[6]), .A1(n3), .B0(b[6]), .B1(n4), .Y(n14) );
  AOI22XL U4 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  AOI22XL U5 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n4), .Y(n15) );
  INVX1 U6 ( .A(n2), .Y(n3) );
  INVX1 U7 ( .A(n1), .Y(n4) );
  INVX1 U8 ( .A(n2), .Y(n1) );
  INVX1 U9 ( .A(sel), .Y(n2) );
  INVX1 U10 ( .A(n6), .Y(out[10]) );
  INVX1 U11 ( .A(n9), .Y(out[1]) );
  AOI22X1 U12 ( .A0(a[1]), .A1(n3), .B0(b[1]), .B1(n2), .Y(n9) );
  INVX1 U13 ( .A(n8), .Y(out[12]) );
  INVX1 U14 ( .A(n7), .Y(out[11]) );
  INVX1 U15 ( .A(n18), .Y(out[9]) );
  INVX1 U16 ( .A(n17), .Y(out[8]) );
  INVX1 U17 ( .A(n15), .Y(out[7]) );
  INVX1 U18 ( .A(n14), .Y(out[6]) );
  INVX1 U19 ( .A(n13), .Y(out[5]) );
  AOI22X1 U20 ( .A0(a[5]), .A1(n3), .B0(b[5]), .B1(n2), .Y(n13) );
  INVX1 U21 ( .A(n12), .Y(out[4]) );
  AOI22X1 U22 ( .A0(a[4]), .A1(n3), .B0(b[4]), .B1(n2), .Y(n12) );
  INVX1 U23 ( .A(n11), .Y(out[3]) );
  AOI22X1 U24 ( .A0(a[3]), .A1(n3), .B0(b[3]), .B1(n4), .Y(n11) );
  INVX1 U25 ( .A(n10), .Y(out[2]) );
  AOI22X1 U26 ( .A0(a[2]), .A1(n3), .B0(b[2]), .B1(n2), .Y(n10) );
  INVX1 U27 ( .A(n5), .Y(out[0]) );
  AOI22X1 U28 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n2), .Y(n5) );
  AOI22X1 U29 ( .A0(a[11]), .A1(n3), .B0(b[11]), .B1(n4), .Y(n7) );
  AOI22XL U30 ( .A0(a[12]), .A1(n3), .B0(b[12]), .B1(n2), .Y(n8) );
endmodule


module mux_13_6 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  AOI22XL U1 ( .A0(a[3]), .A1(n3), .B0(b[3]), .B1(n4), .Y(n11) );
  AOI22XL U2 ( .A0(a[5]), .A1(n3), .B0(b[5]), .B1(n2), .Y(n13) );
  AOI22XL U3 ( .A0(a[12]), .A1(n3), .B0(b[12]), .B1(n2), .Y(n8) );
  AOI22XL U4 ( .A0(a[11]), .A1(n3), .B0(b[11]), .B1(n4), .Y(n7) );
  AOI22XL U5 ( .A0(a[10]), .A1(n3), .B0(b[10]), .B1(n4), .Y(n6) );
  AOI22XL U6 ( .A0(a[6]), .A1(n3), .B0(b[6]), .B1(n4), .Y(n14) );
  AOI22XL U7 ( .A0(a[4]), .A1(n3), .B0(b[4]), .B1(n2), .Y(n12) );
  AOI22XL U8 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n4), .Y(n5) );
  AOI22XL U9 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n17) );
  AOI22XL U10 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n4), .Y(n15) );
  INVX1 U11 ( .A(n2), .Y(n3) );
  INVX1 U12 ( .A(n1), .Y(n4) );
  INVX1 U13 ( .A(n2), .Y(n1) );
  INVX1 U14 ( .A(sel), .Y(n2) );
  INVX1 U15 ( .A(n8), .Y(out[12]) );
  INVX1 U16 ( .A(n7), .Y(out[11]) );
  INVX1 U17 ( .A(n6), .Y(out[10]) );
  INVX1 U18 ( .A(n18), .Y(out[9]) );
  AOI22X1 U19 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  INVX1 U20 ( .A(n17), .Y(out[8]) );
  INVX1 U21 ( .A(n15), .Y(out[7]) );
  INVX1 U22 ( .A(n14), .Y(out[6]) );
  INVX1 U23 ( .A(n13), .Y(out[5]) );
  INVX1 U24 ( .A(n12), .Y(out[4]) );
  INVX1 U25 ( .A(n11), .Y(out[3]) );
  INVX1 U26 ( .A(n10), .Y(out[2]) );
  AOI22X1 U27 ( .A0(a[2]), .A1(n3), .B0(b[2]), .B1(n4), .Y(n10) );
  INVX1 U28 ( .A(n9), .Y(out[1]) );
  AOI22X1 U29 ( .A0(a[1]), .A1(n3), .B0(b[1]), .B1(n2), .Y(n9) );
  INVX1 U30 ( .A(n5), .Y(out[0]) );
endmodule


module mux_13_5 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n3), .Y(n15) );
  AOI22XL U2 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n3), .Y(n7) );
  AOI22XL U3 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n3), .Y(n6) );
  AOI22XL U4 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n1), .Y(n5) );
  AOI22XL U5 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  AOI22XL U6 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n1), .Y(n14) );
  INVX1 U7 ( .A(n1), .Y(n2) );
  INVX1 U8 ( .A(sel), .Y(n3) );
  INVX1 U9 ( .A(sel), .Y(n1) );
  INVX1 U10 ( .A(n7), .Y(out[12]) );
  INVX1 U11 ( .A(n6), .Y(out[11]) );
  INVX1 U12 ( .A(n5), .Y(out[10]) );
  INVX1 U13 ( .A(n17), .Y(out[9]) );
  INVX1 U14 ( .A(n15), .Y(out[8]) );
  INVX1 U15 ( .A(n14), .Y(out[7]) );
  INVX1 U16 ( .A(n13), .Y(out[6]) );
  AOI22X1 U17 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n1), .Y(n13) );
  INVX1 U18 ( .A(n12), .Y(out[5]) );
  AOI22X1 U19 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n3), .Y(n12) );
  INVX1 U20 ( .A(n11), .Y(out[4]) );
  AOI22X1 U21 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n3), .Y(n11) );
  INVX1 U22 ( .A(n10), .Y(out[3]) );
  AOI22X1 U23 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n3), .Y(n10) );
  INVX1 U24 ( .A(n9), .Y(out[2]) );
  AOI22X1 U25 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n1), .Y(n9) );
  INVX1 U26 ( .A(n8), .Y(out[1]) );
  AOI22X1 U27 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n8) );
  INVX1 U28 ( .A(n4), .Y(out[0]) );
  AOI22X1 U29 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n4) );
endmodule


module mux_13_4 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  INVX1 U1 ( .A(sel), .Y(n1) );
  AOI22XL U2 ( .A0(a[7]), .A1(n2), .B0(b[7]), .B1(n3), .Y(n14) );
  AOI22XL U3 ( .A0(a[8]), .A1(n2), .B0(b[8]), .B1(n3), .Y(n15) );
  AOI22XL U4 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  AOI22XL U5 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n1), .Y(n4) );
  AOI22XL U6 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n3), .Y(n10) );
  AOI22XL U7 ( .A0(a[12]), .A1(sel), .B0(b[12]), .B1(n1), .Y(n7) );
  AOI22XL U8 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n13) );
  AOI22XL U9 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n3), .Y(n8) );
  AOI22XL U10 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n3), .Y(n12) );
  AOI22XL U11 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n3), .Y(n6) );
  AOI22XL U12 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n3), .Y(n11) );
  AOI22XL U13 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n3), .Y(n5) );
  INVX1 U14 ( .A(n17), .Y(out[9]) );
  INVX1 U15 ( .A(n15), .Y(out[8]) );
  INVX1 U16 ( .A(n14), .Y(out[7]) );
  BUFX3 U17 ( .A(n1), .Y(n3) );
  BUFX3 U18 ( .A(sel), .Y(n2) );
  INVX1 U19 ( .A(n13), .Y(out[6]) );
  INVX1 U20 ( .A(n10), .Y(out[3]) );
  INVX1 U21 ( .A(n7), .Y(out[12]) );
  INVX1 U22 ( .A(n4), .Y(out[0]) );
  INVX1 U23 ( .A(n12), .Y(out[5]) );
  INVX1 U24 ( .A(n9), .Y(out[2]) );
  AOI22X1 U25 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n1), .Y(n9) );
  INVX1 U26 ( .A(n6), .Y(out[11]) );
  INVX1 U27 ( .A(n11), .Y(out[4]) );
  INVX1 U28 ( .A(n8), .Y(out[1]) );
  INVX1 U29 ( .A(n5), .Y(out[10]) );
endmodule


module mux_13_3 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n3), .Y(n9) );
  AOI22XL U2 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n3), .Y(n8) );
  AOI22XL U3 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n3), .Y(n7) );
  AOI22XL U4 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n2), .Y(n6) );
  AOI22XL U5 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n5) );
  AOI22XL U6 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n2), .Y(n13) );
  AOI22XL U7 ( .A0(a[5]), .A1(sel), .B0(b[5]), .B1(n2), .Y(n12) );
  AOI22XL U8 ( .A0(a[4]), .A1(sel), .B0(b[4]), .B1(n3), .Y(n11) );
  AOI22XL U9 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n2), .Y(n10) );
  AOI22XL U10 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n4) );
  AOI22XL U11 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n3), .Y(n17) );
  AOI22XL U12 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n2), .Y(n15) );
  AOI22XL U13 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n2), .Y(n14) );
  INVX1 U14 ( .A(n1), .Y(n3) );
  INVX1 U15 ( .A(n2), .Y(n1) );
  INVX1 U16 ( .A(n7), .Y(out[12]) );
  INVX1 U17 ( .A(n6), .Y(out[11]) );
  INVX1 U18 ( .A(n5), .Y(out[10]) );
  INVX1 U19 ( .A(n17), .Y(out[9]) );
  INVX1 U20 ( .A(n15), .Y(out[8]) );
  INVX1 U21 ( .A(n14), .Y(out[7]) );
  INVX1 U22 ( .A(n13), .Y(out[6]) );
  INVX1 U23 ( .A(n12), .Y(out[5]) );
  INVX1 U24 ( .A(n11), .Y(out[4]) );
  INVX1 U25 ( .A(n10), .Y(out[3]) );
  INVX1 U26 ( .A(n9), .Y(out[2]) );
  INVX1 U27 ( .A(n8), .Y(out[1]) );
  INVX1 U28 ( .A(n4), .Y(out[0]) );
  INVX1 U29 ( .A(sel), .Y(n2) );
endmodule


module mux_13_2 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n5) );
  AOI22XL U2 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n3), .Y(n13) );
  AOI22XL U3 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n12) );
  AOI22XL U4 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n17) );
  AOI22XL U5 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n2), .Y(n15) );
  AOI22XL U6 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n2), .Y(n14) );
  INVX1 U7 ( .A(n3), .Y(n1) );
  INVX1 U8 ( .A(sel), .Y(n2) );
  INVX1 U9 ( .A(sel), .Y(n3) );
  INVX1 U10 ( .A(n5), .Y(out[10]) );
  INVX1 U11 ( .A(n8), .Y(out[1]) );
  AOI22X1 U12 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n3), .Y(n8) );
  INVX1 U13 ( .A(n7), .Y(out[12]) );
  INVX1 U14 ( .A(n6), .Y(out[11]) );
  INVX1 U15 ( .A(n17), .Y(out[9]) );
  INVX1 U16 ( .A(n15), .Y(out[8]) );
  INVX1 U17 ( .A(n14), .Y(out[7]) );
  INVX1 U18 ( .A(n13), .Y(out[6]) );
  INVX1 U19 ( .A(n12), .Y(out[5]) );
  INVX1 U20 ( .A(n11), .Y(out[4]) );
  AOI22X1 U21 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n2), .Y(n11) );
  INVX1 U22 ( .A(n10), .Y(out[3]) );
  AOI22X1 U23 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n2), .Y(n10) );
  INVX1 U24 ( .A(n9), .Y(out[2]) );
  AOI22X1 U25 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n9) );
  INVX1 U26 ( .A(n4), .Y(out[0]) );
  AOI22X1 U27 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n4) );
  AOI22XL U28 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n3), .Y(n7) );
  AOI22XL U29 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n2), .Y(n6) );
endmodule


module mux_13_1 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n20, n21, n22;

  AOI22XL U1 ( .A0(a[6]), .A1(n3), .B0(b[6]), .B1(n4), .Y(n17) );
  AOI22XL U2 ( .A0(a[12]), .A1(n3), .B0(b[12]), .B1(n6), .Y(n10) );
  AOI22XL U3 ( .A0(a[11]), .A1(n3), .B0(b[11]), .B1(n6), .Y(n9) );
  AOI22XL U4 ( .A0(a[10]), .A1(n3), .B0(b[10]), .B1(n6), .Y(n8) );
  AOI22XL U5 ( .A0(a[1]), .A1(n3), .B0(b[1]), .B1(n5), .Y(n11) );
  AOI22XL U6 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n2), .Y(n7) );
  AOI22XL U7 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n5), .Y(n21) );
  AOI22XL U8 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n4), .Y(n20) );
  INVX1 U9 ( .A(n2), .Y(n3) );
  INVX1 U10 ( .A(n1), .Y(n6) );
  INVX1 U11 ( .A(n1), .Y(n4) );
  INVX1 U12 ( .A(n1), .Y(n5) );
  INVX1 U13 ( .A(n2), .Y(n1) );
  INVX1 U14 ( .A(sel), .Y(n2) );
  INVX1 U15 ( .A(n10), .Y(out[12]) );
  INVX1 U16 ( .A(n9), .Y(out[11]) );
  INVX1 U17 ( .A(n8), .Y(out[10]) );
  INVX1 U18 ( .A(n22), .Y(out[9]) );
  AOI22X1 U19 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n22) );
  INVX1 U20 ( .A(n21), .Y(out[8]) );
  INVX1 U21 ( .A(n20), .Y(out[7]) );
  INVX1 U22 ( .A(n17), .Y(out[6]) );
  INVX1 U23 ( .A(n15), .Y(out[5]) );
  AOI22X1 U24 ( .A0(a[5]), .A1(n3), .B0(b[5]), .B1(n4), .Y(n15) );
  INVX1 U25 ( .A(n14), .Y(out[4]) );
  AOI22X1 U26 ( .A0(a[4]), .A1(n3), .B0(b[4]), .B1(n4), .Y(n14) );
  INVX1 U27 ( .A(n13), .Y(out[3]) );
  AOI22X1 U28 ( .A0(a[3]), .A1(n3), .B0(b[3]), .B1(n5), .Y(n13) );
  INVX1 U29 ( .A(n12), .Y(out[2]) );
  AOI22X1 U30 ( .A0(a[2]), .A1(n3), .B0(b[2]), .B1(n5), .Y(n12) );
  INVX1 U31 ( .A(n11), .Y(out[1]) );
  INVX1 U32 ( .A(n7), .Y(out[0]) );
endmodule


module mux_13_0 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  AOI22XL U1 ( .A0(a[3]), .A1(n2), .B0(b[3]), .B1(n3), .Y(n10) );
  AOI22XL U2 ( .A0(a[2]), .A1(n2), .B0(b[2]), .B1(n1), .Y(n9) );
  AOI22XL U3 ( .A0(a[12]), .A1(n2), .B0(b[12]), .B1(n3), .Y(n7) );
  AOI22XL U4 ( .A0(a[11]), .A1(n2), .B0(b[11]), .B1(n3), .Y(n6) );
  AOI22XL U5 ( .A0(a[10]), .A1(n2), .B0(b[10]), .B1(n1), .Y(n5) );
  AOI22XL U6 ( .A0(a[6]), .A1(n2), .B0(b[6]), .B1(n3), .Y(n13) );
  AOI22XL U7 ( .A0(a[5]), .A1(n2), .B0(b[5]), .B1(n3), .Y(n12) );
  AOI22XL U8 ( .A0(a[4]), .A1(n2), .B0(b[4]), .B1(n3), .Y(n11) );
  AOI22XL U9 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n1), .Y(n17) );
  AOI22XL U10 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n1), .Y(n15) );
  AOI22XL U11 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n3), .Y(n14) );
  INVX1 U12 ( .A(n1), .Y(n2) );
  INVX1 U13 ( .A(sel), .Y(n3) );
  INVX1 U14 ( .A(sel), .Y(n1) );
  INVX1 U15 ( .A(n7), .Y(out[12]) );
  INVX1 U16 ( .A(n6), .Y(out[11]) );
  INVX1 U17 ( .A(n5), .Y(out[10]) );
  INVX1 U18 ( .A(n17), .Y(out[9]) );
  INVX1 U19 ( .A(n15), .Y(out[8]) );
  INVX1 U20 ( .A(n14), .Y(out[7]) );
  INVX1 U21 ( .A(n13), .Y(out[6]) );
  INVX1 U22 ( .A(n12), .Y(out[5]) );
  INVX1 U23 ( .A(n11), .Y(out[4]) );
  INVX1 U24 ( .A(n10), .Y(out[3]) );
  INVX1 U25 ( .A(n9), .Y(out[2]) );
  INVX1 U26 ( .A(n8), .Y(out[1]) );
  AOI22X1 U27 ( .A0(a[1]), .A1(n2), .B0(b[1]), .B1(n1), .Y(n8) );
  INVX1 U28 ( .A(n4), .Y(out[0]) );
  AOI22X1 U29 ( .A0(a[0]), .A1(n2), .B0(b[0]), .B1(n3), .Y(n4) );
endmodule


module mux_5_2to1_0 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7;

  INVX1 U1 ( .A(n2), .Y(n1) );
  INVX1 U2 ( .A(sel), .Y(n2) );
  INVX1 U3 ( .A(n6), .Y(out[3]) );
  AOI22X1 U4 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n2), .Y(n6) );
  INVX1 U5 ( .A(n4), .Y(out[1]) );
  AOI22X1 U6 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n4) );
  INVX1 U7 ( .A(n3), .Y(out[0]) );
  AOI22X1 U8 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n3) );
  INVX1 U9 ( .A(n5), .Y(out[2]) );
  AOI22X1 U10 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n5) );
  INVX1 U11 ( .A(n7), .Y(out[4]) );
  AOI22X1 U12 ( .A0(n1), .A1(a[4]), .B0(b[4]), .B1(n2), .Y(n7) );
endmodule


module mux_5_22 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n4), .Y(out[3]) );
  AOI22X1 U3 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U4 ( .A(n3), .Y(out[2]) );
  AOI22X1 U5 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U6 ( .A(n2), .Y(out[1]) );
  AOI22X1 U7 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U8 ( .A(n1), .Y(out[0]) );
  AOI22X1 U9 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U10 ( .A(n6), .Y(out[4]) );
  AOI22X1 U11 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
endmodule


module mux_5_21 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
  INVX1 U4 ( .A(n4), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U6 ( .A(n1), .Y(out[0]) );
  AOI22X1 U7 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U8 ( .A(n2), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U10 ( .A(n3), .Y(out[2]) );
  AOI22X1 U11 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
endmodule


module mux_5_20 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
  INVX1 U4 ( .A(n4), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U6 ( .A(n3), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U8 ( .A(n2), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U10 ( .A(n1), .Y(out[0]) );
  AOI22X1 U11 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
endmodule


module mux_5_19 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7;

  INVX1 U1 ( .A(n2), .Y(n1) );
  INVX1 U2 ( .A(sel), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(out[0]) );
  AOI22X1 U4 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n3) );
  INVX1 U5 ( .A(n4), .Y(out[1]) );
  AOI22X1 U6 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(out[2]) );
  AOI22X1 U8 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n5) );
  INVX1 U9 ( .A(n6), .Y(out[3]) );
  AOI22X1 U10 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n2), .Y(n6) );
  INVX1 U11 ( .A(n7), .Y(out[4]) );
  AOI22X1 U12 ( .A0(n1), .A1(a[4]), .B0(b[4]), .B1(n2), .Y(n7) );
endmodule


module mux_5_18 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n1) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n1), .Y(n6) );
  INVX1 U4 ( .A(n5), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n1), .Y(n5) );
  INVX1 U6 ( .A(n4), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n1), .Y(n4) );
  INVX1 U8 ( .A(n3), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n1), .Y(n3) );
  INVX1 U10 ( .A(n2), .Y(out[0]) );
  AOI22X1 U11 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n1), .Y(n2) );
endmodule


module mux_5_17 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n1), .Y(out[0]) );
  AOI22X1 U3 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U4 ( .A(n2), .Y(out[1]) );
  AOI22X1 U5 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U6 ( .A(n3), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U8 ( .A(n4), .Y(out[3]) );
  AOI22X1 U9 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U10 ( .A(n6), .Y(out[4]) );
  AOI22X1 U11 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
endmodule


module mux_5_16 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n4), .Y(out[3]) );
  AOI22X1 U3 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U4 ( .A(n3), .Y(out[2]) );
  AOI22X1 U5 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U6 ( .A(n2), .Y(out[1]) );
  AOI22X1 U7 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U8 ( .A(n1), .Y(out[0]) );
  AOI22X1 U9 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U10 ( .A(n6), .Y(out[4]) );
  AOI22X1 U11 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
endmodule


module mux_5_15 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
  INVX1 U4 ( .A(n4), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U6 ( .A(n1), .Y(out[0]) );
  AOI22X1 U7 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U8 ( .A(n2), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U10 ( .A(n3), .Y(out[2]) );
  AOI22X1 U11 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
endmodule


module mux_5_14 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
  INVX1 U4 ( .A(n4), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U6 ( .A(n3), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U8 ( .A(n2), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U10 ( .A(n1), .Y(out[0]) );
  AOI22X1 U11 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
endmodule


module mux_5_13 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7;

  INVX1 U1 ( .A(n2), .Y(n1) );
  INVX1 U2 ( .A(sel), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(out[0]) );
  AOI22X1 U4 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n3) );
  INVX1 U5 ( .A(n4), .Y(out[1]) );
  AOI22X1 U6 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(out[2]) );
  AOI22X1 U8 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n5) );
  INVX1 U9 ( .A(n6), .Y(out[3]) );
  AOI22X1 U10 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n2), .Y(n6) );
  INVX1 U11 ( .A(n7), .Y(out[4]) );
  AOI22X1 U12 ( .A0(n1), .A1(a[4]), .B0(b[4]), .B1(n2), .Y(n7) );
endmodule


module mux_5_12 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n1) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n1), .Y(n6) );
  INVX1 U4 ( .A(n5), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n1), .Y(n5) );
  INVX1 U6 ( .A(n4), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n1), .Y(n4) );
  INVX1 U8 ( .A(n3), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n1), .Y(n3) );
  INVX1 U10 ( .A(n2), .Y(out[0]) );
  AOI22X1 U11 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n1), .Y(n2) );
endmodule


module mux_5_11 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n1), .Y(out[0]) );
  AOI22X1 U3 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U4 ( .A(n2), .Y(out[1]) );
  AOI22X1 U5 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U6 ( .A(n3), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U8 ( .A(n4), .Y(out[3]) );
  AOI22X1 U9 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U10 ( .A(n6), .Y(out[4]) );
  AOI22X1 U11 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
endmodule


module mux_5_10 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n4), .Y(out[3]) );
  AOI22X1 U3 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U4 ( .A(n3), .Y(out[2]) );
  AOI22X1 U5 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U6 ( .A(n2), .Y(out[1]) );
  AOI22X1 U7 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U8 ( .A(n1), .Y(out[0]) );
  AOI22X1 U9 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U10 ( .A(n6), .Y(out[4]) );
  AOI22X1 U11 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
endmodule


module mux_5_9 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
  INVX1 U4 ( .A(n4), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U6 ( .A(n1), .Y(out[0]) );
  AOI22X1 U7 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U8 ( .A(n2), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U10 ( .A(n3), .Y(out[2]) );
  AOI22X1 U11 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
endmodule


module mux_5_8 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
  INVX1 U4 ( .A(n4), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U6 ( .A(n3), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U8 ( .A(n2), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U10 ( .A(n1), .Y(out[0]) );
  AOI22X1 U11 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
endmodule


module mux_5_7 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7;

  INVX1 U1 ( .A(n2), .Y(n1) );
  INVX1 U2 ( .A(sel), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(out[0]) );
  AOI22X1 U4 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n3) );
  INVX1 U5 ( .A(n4), .Y(out[1]) );
  AOI22X1 U6 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(out[2]) );
  AOI22X1 U8 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n5) );
  INVX1 U9 ( .A(n6), .Y(out[3]) );
  AOI22X1 U10 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n2), .Y(n6) );
  INVX1 U11 ( .A(n7), .Y(out[4]) );
  AOI22X1 U12 ( .A0(n1), .A1(a[4]), .B0(b[4]), .B1(n2), .Y(n7) );
endmodule


module mux_5_6 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n1) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n1), .Y(n6) );
  INVX1 U4 ( .A(n5), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n1), .Y(n5) );
  INVX1 U6 ( .A(n4), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n1), .Y(n4) );
  INVX1 U8 ( .A(n3), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n1), .Y(n3) );
  INVX1 U10 ( .A(n2), .Y(out[0]) );
  AOI22X1 U11 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n1), .Y(n2) );
endmodule


module mux_5_5 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n1), .Y(out[0]) );
  AOI22X1 U3 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U4 ( .A(n2), .Y(out[1]) );
  AOI22X1 U5 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U6 ( .A(n3), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U8 ( .A(n4), .Y(out[3]) );
  AOI22X1 U9 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U10 ( .A(n6), .Y(out[4]) );
  AOI22X1 U11 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
endmodule


module mux_5_4 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n4), .Y(out[3]) );
  AOI22X1 U3 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U4 ( .A(n3), .Y(out[2]) );
  AOI22X1 U5 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U6 ( .A(n2), .Y(out[1]) );
  AOI22X1 U7 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U8 ( .A(n1), .Y(out[0]) );
  AOI22X1 U9 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U10 ( .A(n6), .Y(out[4]) );
  AOI22X1 U11 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
endmodule


module mux_5_3 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
  INVX1 U4 ( .A(n4), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U6 ( .A(n1), .Y(out[0]) );
  AOI22X1 U7 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
  INVX1 U8 ( .A(n2), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U10 ( .A(n3), .Y(out[2]) );
  AOI22X1 U11 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
endmodule


module mux_5_2 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n5) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n5), .Y(n6) );
  INVX1 U4 ( .A(n4), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n5), .Y(n4) );
  INVX1 U6 ( .A(n3), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n5), .Y(n3) );
  INVX1 U8 ( .A(n2), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n5), .Y(n2) );
  INVX1 U10 ( .A(n1), .Y(out[0]) );
  AOI22X1 U11 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n5), .Y(n1) );
endmodule


module mux_5_1 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7;

  INVX1 U1 ( .A(n2), .Y(n1) );
  INVX1 U2 ( .A(sel), .Y(n2) );
  INVX1 U3 ( .A(n3), .Y(out[0]) );
  AOI22X1 U4 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n3) );
  INVX1 U5 ( .A(n4), .Y(out[1]) );
  AOI22X1 U6 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n4) );
  INVX1 U7 ( .A(n5), .Y(out[2]) );
  AOI22X1 U8 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n5) );
  INVX1 U9 ( .A(n6), .Y(out[3]) );
  AOI22X1 U10 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n2), .Y(n6) );
  INVX1 U11 ( .A(n7), .Y(out[4]) );
  AOI22X1 U12 ( .A0(n1), .A1(a[4]), .B0(b[4]), .B1(n2), .Y(n7) );
endmodule


module mux_5_0 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6;

  INVX1 U1 ( .A(sel), .Y(n1) );
  INVX1 U2 ( .A(n6), .Y(out[4]) );
  AOI22X1 U3 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n1), .Y(n6) );
  INVX1 U4 ( .A(n5), .Y(out[3]) );
  AOI22X1 U5 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n1), .Y(n5) );
  INVX1 U6 ( .A(n4), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n1), .Y(n4) );
  INVX1 U8 ( .A(n3), .Y(out[1]) );
  AOI22X1 U9 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n1), .Y(n3) );
  INVX1 U10 ( .A(n2), .Y(out[0]) );
  AOI22X1 U11 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n1), .Y(n2) );
endmodule


module mux_1_2to1_0 ( a, b, sel, out );
  input a, b, sel;
  output out;
  wire   n1;

  OAI2BB2X1 U1 ( .B0(n1), .B1(sel), .A0N(sel), .A1N(a), .Y(out) );
  INVX1 U2 ( .A(b), .Y(n1) );
endmodule


module mux13_13_7 ( a, b, sel, enable, out, clk, reset );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel, enable, clk, reset;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N83,
         n14, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42;

  EDFFX1 \out_reg[11]  ( .D(N28), .E(N83), .CK(clk), .Q(out[11]) );
  EDFFX1 \out_reg[9]  ( .D(N26), .E(N83), .CK(clk), .Q(out[9]) );
  EDFFX1 \out_reg[8]  ( .D(N25), .E(N83), .CK(clk), .Q(out[8]) );
  EDFFX1 \out_reg[7]  ( .D(N24), .E(N83), .CK(clk), .Q(out[7]) );
  EDFFX1 \out_reg[6]  ( .D(N23), .E(N83), .CK(clk), .Q(out[6]) );
  EDFFX1 \out_reg[5]  ( .D(N22), .E(N83), .CK(clk), .Q(out[5]) );
  EDFFX1 \out_reg[4]  ( .D(N21), .E(N83), .CK(clk), .Q(out[4]) );
  EDFFX1 \out_reg[0]  ( .D(N17), .E(N83), .CK(clk), .Q(out[0]) );
  EDFFX1 \out_reg[2]  ( .D(N19), .E(N83), .CK(clk), .Q(out[2]) );
  EDFFX1 \out_reg[3]  ( .D(N20), .E(N83), .CK(clk), .Q(out[3]) );
  EDFFX1 \out_reg[1]  ( .D(N18), .E(N83), .CK(clk), .Q(out[1]) );
  EDFFX1 \out_reg[10]  ( .D(N27), .E(N83), .CK(clk), .Q(out[10]) );
  EDFFX1 \out_reg[12]  ( .D(N29), .E(N83), .CK(clk), .Q(out[12]) );
  AOI22XL U3 ( .A0(b[10]), .A1(n41), .B0(a[10]), .B1(n40), .Y(n38) );
  AOI22XL U4 ( .A0(b[0]), .A1(n41), .B0(a[0]), .B1(n40), .Y(n14) );
  INVX1 U5 ( .A(n29), .Y(N18) );
  AOI22X1 U6 ( .A0(b[1]), .A1(n41), .B0(a[1]), .B1(n40), .Y(n29) );
  INVX1 U7 ( .A(n33), .Y(N22) );
  AOI22X1 U8 ( .A0(b[5]), .A1(n41), .B0(a[5]), .B1(n40), .Y(n33) );
  INVX1 U9 ( .A(n32), .Y(N21) );
  AOI22X1 U10 ( .A0(b[4]), .A1(n41), .B0(a[4]), .B1(n40), .Y(n32) );
  INVX1 U11 ( .A(n31), .Y(N20) );
  AOI22X1 U12 ( .A0(b[3]), .A1(n41), .B0(a[3]), .B1(n40), .Y(n31) );
  INVX1 U13 ( .A(n39), .Y(N28) );
  AOI22X1 U14 ( .A0(b[11]), .A1(n41), .B0(a[11]), .B1(n40), .Y(n39) );
  NAND2BX1 U15 ( .AN(enable), .B(reset), .Y(N83) );
  INVX1 U16 ( .A(n34), .Y(N23) );
  AOI22X1 U17 ( .A0(b[6]), .A1(n41), .B0(a[6]), .B1(n40), .Y(n34) );
  INVX1 U18 ( .A(n35), .Y(N24) );
  AOI22X1 U19 ( .A0(b[7]), .A1(n41), .B0(a[7]), .B1(n40), .Y(n35) );
  INVX1 U20 ( .A(n42), .Y(N29) );
  AOI22X1 U21 ( .A0(b[12]), .A1(n41), .B0(a[12]), .B1(n40), .Y(n42) );
  INVX1 U22 ( .A(n14), .Y(N17) );
  INVX1 U23 ( .A(n30), .Y(N19) );
  AOI22X1 U24 ( .A0(b[2]), .A1(n41), .B0(a[2]), .B1(n40), .Y(n30) );
  INVX1 U25 ( .A(n36), .Y(N25) );
  AOI22X1 U26 ( .A0(b[8]), .A1(n41), .B0(a[8]), .B1(n40), .Y(n36) );
  INVX1 U27 ( .A(n37), .Y(N26) );
  AOI22X1 U28 ( .A0(b[9]), .A1(n41), .B0(a[9]), .B1(n40), .Y(n37) );
  INVX1 U29 ( .A(n38), .Y(N27) );
  NOR2BX1 U30 ( .AN(reset), .B(sel), .Y(n41) );
  AND2X2 U31 ( .A(sel), .B(reset), .Y(n40) );
endmodule


module mux13_13_6 ( a, b, sel, enable, out, clk, reset );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel, enable, clk, reset;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N83,
         n5, n12, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42;

  EDFFX4 \out_reg[12]  ( .D(N29), .E(N83), .CK(clk), .Q(out[12]) );
  EDFFX4 \out_reg[11]  ( .D(N28), .E(N83), .CK(clk), .Q(out[11]) );
  EDFFX4 \out_reg[9]  ( .D(N26), .E(N83), .CK(clk), .Q(out[9]) );
  EDFFX4 \out_reg[7]  ( .D(N24), .E(N83), .CK(clk), .Q(out[7]) );
  EDFFX4 \out_reg[1]  ( .D(N18), .E(N83), .CK(clk), .Q(out[1]) );
  EDFFX4 \out_reg[0]  ( .D(N17), .E(N83), .CK(clk), .Q(out[0]) );
  EDFFX1 \out_reg[5]  ( .D(N22), .E(N83), .CK(clk), .Q(out[5]) );
  EDFFX1 \out_reg[4]  ( .D(N21), .E(N83), .CK(clk), .Q(out[4]) );
  EDFFX1 \out_reg[3]  ( .D(N20), .E(N83), .CK(clk), .Q(out[3]) );
  EDFFX2 \out_reg[6]  ( .D(N23), .E(N83), .CK(clk), .Q(out[6]) );
  MX2X1 \out_reg[2]/U3  ( .A(out[2]), .B(N19), .S0(N83), .Y(n5) );
  DFFHQX2 \out_reg[2]  ( .D(n5), .CK(clk), .Q(out[2]) );
  EDFFX2 \out_reg[8]  ( .D(N25), .E(N83), .CK(clk), .Q(out[8]) );
  EDFFX4 \out_reg[10]  ( .D(N27), .E(N83), .CK(clk), .Q(out[10]) );
  AOI22XL U3 ( .A0(b[6]), .A1(n41), .B0(a[6]), .B1(n40), .Y(n34) );
  AOI22XL U4 ( .A0(b[4]), .A1(n41), .B0(a[4]), .B1(n40), .Y(n32) );
  AOI22XL U5 ( .A0(b[5]), .A1(n41), .B0(a[5]), .B1(n40), .Y(n33) );
  AOI22XL U6 ( .A0(b[7]), .A1(n41), .B0(a[7]), .B1(n40), .Y(n35) );
  AOI22XL U7 ( .A0(b[8]), .A1(n41), .B0(a[8]), .B1(n40), .Y(n36) );
  AOI22XL U8 ( .A0(b[9]), .A1(n41), .B0(a[9]), .B1(n40), .Y(n37) );
  AOI22XL U9 ( .A0(b[11]), .A1(n41), .B0(a[11]), .B1(n40), .Y(n39) );
  INVX1 U10 ( .A(n32), .Y(N21) );
  INVX1 U11 ( .A(n33), .Y(N22) );
  INVX1 U12 ( .A(n34), .Y(N23) );
  INVX1 U13 ( .A(n29), .Y(N18) );
  AOI22X1 U14 ( .A0(b[1]), .A1(n41), .B0(a[1]), .B1(n40), .Y(n29) );
  INVX1 U15 ( .A(n38), .Y(N27) );
  INVX1 U16 ( .A(n12), .Y(N17) );
  AOI22XL U17 ( .A0(b[0]), .A1(n41), .B0(a[0]), .B1(n40), .Y(n12) );
  INVX1 U18 ( .A(n31), .Y(N20) );
  AOI22X1 U19 ( .A0(b[3]), .A1(n41), .B0(a[3]), .B1(n40), .Y(n31) );
  INVX1 U20 ( .A(n35), .Y(N24) );
  INVX1 U21 ( .A(n36), .Y(N25) );
  INVX1 U22 ( .A(n37), .Y(N26) );
  INVX1 U23 ( .A(n39), .Y(N28) );
  INVX1 U24 ( .A(n42), .Y(N29) );
  AOI22X1 U25 ( .A0(b[12]), .A1(n41), .B0(a[12]), .B1(n40), .Y(n42) );
  NOR2BX1 U26 ( .AN(reset), .B(sel), .Y(n41) );
  AND2X2 U27 ( .A(sel), .B(reset), .Y(n40) );
  NAND2BX1 U28 ( .AN(enable), .B(reset), .Y(N83) );
  INVX1 U29 ( .A(n30), .Y(N19) );
  AOI22X1 U30 ( .A0(b[2]), .A1(n41), .B0(a[2]), .B1(n40), .Y(n30) );
  AOI22X1 U31 ( .A0(b[10]), .A1(n41), .B0(a[10]), .B1(n40), .Y(n38) );
endmodule


module mux13_13_5 ( a, b, sel, enable, out, clk, reset );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel, enable, clk, reset;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N83,
         n8, n9, n10, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42;

  EDFFX4 \out_reg[12]  ( .D(N29), .E(N83), .CK(clk), .Q(out[12]) );
  EDFFX4 \out_reg[11]  ( .D(N28), .E(N83), .CK(clk), .Q(out[11]) );
  EDFFX4 \out_reg[10]  ( .D(N27), .E(N83), .CK(clk), .Q(out[10]) );
  EDFFX4 \out_reg[9]  ( .D(N26), .E(N83), .CK(clk), .Q(out[9]) );
  EDFFX4 \out_reg[4]  ( .D(N21), .E(N83), .CK(clk), .Q(out[4]) );
  EDFFX4 \out_reg[3]  ( .D(N20), .E(N83), .CK(clk), .Q(out[3]) );
  EDFFX4 \out_reg[2]  ( .D(N19), .E(N83), .CK(clk), .Q(out[2]) );
  EDFFX4 \out_reg[1]  ( .D(N18), .E(N83), .CK(clk), .Q(out[1]) );
  EDFFX4 \out_reg[0]  ( .D(N17), .E(N83), .CK(clk), .Q(out[0]) );
  MX2X1 \out_reg[7]/U3  ( .A(out[7]), .B(N24), .S0(N83), .Y(n9) );
  DFFHQX4 \out_reg[7]  ( .D(n9), .CK(clk), .Q(out[7]) );
  MX2X1 \out_reg[8]/U3  ( .A(out[8]), .B(N25), .S0(N83), .Y(n8) );
  DFFHQX4 \out_reg[8]  ( .D(n8), .CK(clk), .Q(out[8]) );
  EDFFX2 \out_reg[5]  ( .D(N22), .E(N83), .CK(clk), .Q(out[5]) );
  EDFFX2 \out_reg[6]  ( .D(N23), .E(N83), .CK(clk), .Q(out[6]) );
  AOI22XL U3 ( .A0(b[2]), .A1(n41), .B0(a[2]), .B1(n40), .Y(n30) );
  INVX1 U4 ( .A(n42), .Y(N29) );
  AOI22X1 U5 ( .A0(b[12]), .A1(n41), .B0(a[12]), .B1(n40), .Y(n42) );
  INVX1 U6 ( .A(n38), .Y(N27) );
  AOI22X1 U7 ( .A0(b[10]), .A1(n41), .B0(a[10]), .B1(n40), .Y(n38) );
  INVX1 U8 ( .A(n39), .Y(N28) );
  AOI22X1 U9 ( .A0(b[11]), .A1(n41), .B0(a[11]), .B1(n40), .Y(n39) );
  INVX1 U10 ( .A(n37), .Y(N26) );
  AOI22X1 U11 ( .A0(b[9]), .A1(n41), .B0(a[9]), .B1(n40), .Y(n37) );
  INVX1 U12 ( .A(n10), .Y(N17) );
  AOI22XL U13 ( .A0(b[0]), .A1(n41), .B0(a[0]), .B1(n40), .Y(n10) );
  NAND2BX1 U14 ( .AN(enable), .B(reset), .Y(N83) );
  INVX1 U15 ( .A(n29), .Y(N18) );
  AOI22X1 U16 ( .A0(b[1]), .A1(n41), .B0(a[1]), .B1(n40), .Y(n29) );
  INVX1 U17 ( .A(n30), .Y(N19) );
  INVX1 U18 ( .A(n33), .Y(N22) );
  AOI22X1 U19 ( .A0(b[5]), .A1(n41), .B0(a[5]), .B1(n40), .Y(n33) );
  INVX1 U20 ( .A(n34), .Y(N23) );
  AOI22X1 U21 ( .A0(b[6]), .A1(n41), .B0(a[6]), .B1(n40), .Y(n34) );
  INVX1 U22 ( .A(n36), .Y(N25) );
  AOI22X1 U23 ( .A0(b[8]), .A1(n41), .B0(a[8]), .B1(n40), .Y(n36) );
  INVX1 U24 ( .A(n35), .Y(N24) );
  AOI22X1 U25 ( .A0(b[7]), .A1(n41), .B0(a[7]), .B1(n40), .Y(n35) );
  INVX1 U26 ( .A(n31), .Y(N20) );
  AOI22XL U27 ( .A0(b[3]), .A1(n41), .B0(a[3]), .B1(n40), .Y(n31) );
  INVX1 U28 ( .A(n32), .Y(N21) );
  AOI22X1 U29 ( .A0(b[4]), .A1(n41), .B0(a[4]), .B1(n40), .Y(n32) );
  NOR2BX1 U30 ( .AN(reset), .B(sel), .Y(n41) );
  AND2X2 U31 ( .A(sel), .B(reset), .Y(n40) );
endmodule


module mux13_13_4 ( a, b, sel, enable, out, clk, reset );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel, enable, clk, reset;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N83,
         n9, n10, n13, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42;

  EDFFX4 \out_reg[12]  ( .D(N29), .E(N83), .CK(clk), .Q(out[12]) );
  EDFFX4 \out_reg[10]  ( .D(N27), .E(N83), .CK(clk), .Q(out[10]) );
  EDFFX4 \out_reg[9]  ( .D(N26), .E(N83), .CK(clk), .Q(out[9]) );
  EDFFX4 \out_reg[6]  ( .D(N23), .E(N83), .CK(clk), .Q(out[6]) );
  EDFFX4 \out_reg[5]  ( .D(N22), .E(N83), .CK(clk), .Q(out[5]) );
  EDFFX4 \out_reg[3]  ( .D(N20), .E(N83), .CK(clk), .Q(out[3]) );
  EDFFX4 \out_reg[1]  ( .D(N18), .E(N83), .CK(clk), .Q(out[1]) );
  MX2X1 \out_reg[2]/U3  ( .A(out[2]), .B(N19), .S0(N83), .Y(n10) );
  DFFHQX4 \out_reg[2]  ( .D(n10), .CK(clk), .Q(out[2]) );
  MX2X1 \out_reg[11]/U3  ( .A(out[11]), .B(N28), .S0(N83), .Y(n9) );
  DFFHQX4 \out_reg[11]  ( .D(n9), .CK(clk), .Q(out[11]) );
  EDFFX1 \out_reg[8]  ( .D(N25), .E(N83), .CK(clk), .Q(out[8]) );
  EDFFX1 \out_reg[0]  ( .D(N17), .E(N83), .CK(clk), .Q(out[0]) );
  EDFFX1 \out_reg[4]  ( .D(N21), .E(N83), .CK(clk), .Q(out[4]) );
  EDFFX2 \out_reg[7]  ( .D(N24), .E(N83), .CK(clk), .Q(out[7]) );
  AOI22XL U3 ( .A0(b[1]), .A1(n41), .B0(a[1]), .B1(n40), .Y(n29) );
  AOI22XL U4 ( .A0(b[2]), .A1(n41), .B0(a[2]), .B1(n40), .Y(n30) );
  AOI22XL U5 ( .A0(b[8]), .A1(n41), .B0(a[8]), .B1(n40), .Y(n36) );
  INVX1 U6 ( .A(n29), .Y(N18) );
  INVX1 U7 ( .A(n31), .Y(N20) );
  AOI22X1 U8 ( .A0(b[3]), .A1(n41), .B0(a[3]), .B1(n40), .Y(n31) );
  INVX1 U9 ( .A(n39), .Y(N28) );
  INVX1 U10 ( .A(n30), .Y(N19) );
  INVX1 U11 ( .A(n13), .Y(N17) );
  AOI22X1 U12 ( .A0(b[0]), .A1(n41), .B0(a[0]), .B1(n40), .Y(n13) );
  INVX1 U13 ( .A(n38), .Y(N27) );
  AOI22X1 U14 ( .A0(b[10]), .A1(n41), .B0(a[10]), .B1(n40), .Y(n38) );
  INVX1 U15 ( .A(n42), .Y(N29) );
  AOI22X1 U16 ( .A0(b[12]), .A1(n41), .B0(a[12]), .B1(n40), .Y(n42) );
  NOR2BX1 U17 ( .AN(reset), .B(sel), .Y(n41) );
  AND2X2 U18 ( .A(sel), .B(reset), .Y(n40) );
  NAND2BX1 U19 ( .AN(enable), .B(reset), .Y(N83) );
  INVX1 U20 ( .A(n32), .Y(N21) );
  AOI22X1 U21 ( .A0(b[4]), .A1(n41), .B0(a[4]), .B1(n40), .Y(n32) );
  INVX1 U22 ( .A(n33), .Y(N22) );
  AOI22X1 U23 ( .A0(b[5]), .A1(n41), .B0(a[5]), .B1(n40), .Y(n33) );
  INVX1 U24 ( .A(n34), .Y(N23) );
  AOI22X1 U25 ( .A0(b[6]), .A1(n41), .B0(a[6]), .B1(n40), .Y(n34) );
  INVX1 U26 ( .A(n35), .Y(N24) );
  AOI22X1 U27 ( .A0(b[7]), .A1(n41), .B0(a[7]), .B1(n40), .Y(n35) );
  INVX1 U28 ( .A(n36), .Y(N25) );
  INVX1 U29 ( .A(n37), .Y(N26) );
  AOI22X1 U30 ( .A0(b[9]), .A1(n41), .B0(a[9]), .B1(n40), .Y(n37) );
  AOI22XL U31 ( .A0(b[11]), .A1(n41), .B0(a[11]), .B1(n40), .Y(n39) );
endmodule


module mux13_13_3 ( a, b, sel, enable, out, clk, reset );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel, enable, clk, reset;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N83,
         n13, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42;

  EDFFX4 \out_reg[12]  ( .D(N29), .E(N83), .CK(clk), .Q(out[12]) );
  EDFFX4 \out_reg[10]  ( .D(N27), .E(N83), .CK(clk), .Q(out[10]) );
  EDFFX4 \out_reg[9]  ( .D(N26), .E(N83), .CK(clk), .Q(out[9]) );
  EDFFX4 \out_reg[8]  ( .D(N25), .E(N83), .CK(clk), .Q(out[8]) );
  EDFFX4 \out_reg[7]  ( .D(N24), .E(N83), .CK(clk), .Q(out[7]) );
  EDFFX4 \out_reg[6]  ( .D(N23), .E(N83), .CK(clk), .Q(out[6]) );
  EDFFX4 \out_reg[5]  ( .D(N22), .E(N83), .CK(clk), .Q(out[5]) );
  EDFFX4 \out_reg[2]  ( .D(N19), .E(N83), .CK(clk), .Q(out[2]) );
  EDFFX4 \out_reg[0]  ( .D(N17), .E(N83), .CK(clk), .Q(out[0]) );
  EDFFX4 \out_reg[1]  ( .D(N18), .E(N83), .CK(clk), .Q(out[1]) );
  EDFFX2 \out_reg[11]  ( .D(N28), .E(N83), .CK(clk), .Q(out[11]) );
  EDFFX2 \out_reg[3]  ( .D(N20), .E(N83), .CK(clk), .Q(out[3]) );
  EDFFX2 \out_reg[4]  ( .D(N21), .E(N83), .CK(clk), .Q(out[4]) );
  AOI22XL U3 ( .A0(b[12]), .A1(n41), .B0(a[12]), .B1(n40), .Y(n42) );
  AOI22XL U4 ( .A0(b[3]), .A1(n41), .B0(a[3]), .B1(n40), .Y(n31) );
  INVX1 U5 ( .A(n35), .Y(N24) );
  AOI22X1 U6 ( .A0(b[7]), .A1(n41), .B0(a[7]), .B1(n40), .Y(n35) );
  INVX1 U7 ( .A(n37), .Y(N26) );
  AOI22X1 U8 ( .A0(b[9]), .A1(n41), .B0(a[9]), .B1(n40), .Y(n37) );
  INVX1 U9 ( .A(n42), .Y(N29) );
  INVX1 U10 ( .A(n13), .Y(N17) );
  AOI22X1 U11 ( .A0(b[0]), .A1(n41), .B0(a[0]), .B1(n40), .Y(n13) );
  INVX1 U12 ( .A(n31), .Y(N20) );
  INVX1 U13 ( .A(n39), .Y(N28) );
  AOI22X1 U14 ( .A0(b[11]), .A1(n41), .B0(a[11]), .B1(n40), .Y(n39) );
  NOR2BX1 U15 ( .AN(reset), .B(sel), .Y(n41) );
  AND2X2 U16 ( .A(sel), .B(reset), .Y(n40) );
  NAND2BX1 U17 ( .AN(enable), .B(reset), .Y(N83) );
  INVX1 U18 ( .A(n29), .Y(N18) );
  AOI22X1 U19 ( .A0(b[1]), .A1(n41), .B0(a[1]), .B1(n40), .Y(n29) );
  INVX1 U20 ( .A(n32), .Y(N21) );
  AOI22X1 U21 ( .A0(b[4]), .A1(n41), .B0(a[4]), .B1(n40), .Y(n32) );
  INVX1 U22 ( .A(n34), .Y(N23) );
  AOI22XL U23 ( .A0(b[6]), .A1(n41), .B0(a[6]), .B1(n40), .Y(n34) );
  INVX1 U24 ( .A(n33), .Y(N22) );
  AOI22X1 U25 ( .A0(b[5]), .A1(n41), .B0(a[5]), .B1(n40), .Y(n33) );
  INVX1 U26 ( .A(n30), .Y(N19) );
  AOI22X1 U27 ( .A0(b[2]), .A1(n41), .B0(a[2]), .B1(n40), .Y(n30) );
  INVX1 U28 ( .A(n36), .Y(N25) );
  AOI22X1 U29 ( .A0(b[8]), .A1(n41), .B0(a[8]), .B1(n40), .Y(n36) );
  INVX1 U30 ( .A(n38), .Y(N27) );
  AOI22X1 U31 ( .A0(b[10]), .A1(n41), .B0(a[10]), .B1(n40), .Y(n38) );
endmodule


module mux13_13_2 ( a, b, sel, enable, out, clk, reset );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel, enable, clk, reset;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N83,
         n14, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42;

  EDFFX4 \out_reg[11]  ( .D(N28), .E(N83), .CK(clk), .Q(out[11]) );
  EDFFX4 \out_reg[10]  ( .D(N27), .E(N83), .CK(clk), .Q(out[10]) );
  EDFFX4 \out_reg[9]  ( .D(N26), .E(N83), .CK(clk), .Q(out[9]) );
  EDFFX4 \out_reg[8]  ( .D(N25), .E(N83), .CK(clk), .Q(out[8]) );
  EDFFX4 \out_reg[5]  ( .D(N22), .E(N83), .CK(clk), .Q(out[5]) );
  EDFFX1 \out_reg[1]  ( .D(N18), .E(N83), .CK(clk), .Q(out[1]) );
  EDFFX4 \out_reg[12]  ( .D(N29), .E(N83), .CK(clk), .Q(out[12]) );
  EDFFX2 \out_reg[2]  ( .D(N19), .E(N83), .CK(clk), .Q(out[2]) );
  EDFFX2 \out_reg[3]  ( .D(N20), .E(N83), .CK(clk), .Q(out[3]) );
  EDFFX2 \out_reg[4]  ( .D(N21), .E(N83), .CK(clk), .Q(out[4]) );
  EDFFX2 \out_reg[7]  ( .D(N24), .E(N83), .CK(clk), .Q(out[7]) );
  EDFFX2 \out_reg[0]  ( .D(N17), .E(N83), .CK(clk), .Q(out[0]) );
  EDFFX2 \out_reg[6]  ( .D(N23), .E(N83), .CK(clk), .Q(out[6]) );
  AOI22XL U3 ( .A0(b[7]), .A1(n41), .B0(a[7]), .B1(n40), .Y(n35) );
  AOI22XL U4 ( .A0(b[2]), .A1(n41), .B0(a[2]), .B1(n40), .Y(n30) );
  INVX1 U5 ( .A(n14), .Y(N17) );
  AOI22X1 U6 ( .A0(b[0]), .A1(n41), .B0(a[0]), .B1(n40), .Y(n14) );
  INVX1 U7 ( .A(n33), .Y(N22) );
  AOI22X1 U8 ( .A0(b[5]), .A1(n41), .B0(a[5]), .B1(n40), .Y(n33) );
  INVX1 U9 ( .A(n37), .Y(N26) );
  AOI22X1 U10 ( .A0(b[9]), .A1(n41), .B0(a[9]), .B1(n40), .Y(n37) );
  INVX1 U11 ( .A(n31), .Y(N20) );
  NOR2BX1 U12 ( .AN(reset), .B(sel), .Y(n41) );
  AND2X2 U13 ( .A(sel), .B(reset), .Y(n40) );
  NAND2BX1 U14 ( .AN(enable), .B(reset), .Y(N83) );
  INVX1 U15 ( .A(n39), .Y(N28) );
  AOI22X1 U16 ( .A0(b[11]), .A1(n41), .B0(a[11]), .B1(n40), .Y(n39) );
  INVX1 U17 ( .A(n32), .Y(N21) );
  AOI22X1 U18 ( .A0(b[4]), .A1(n41), .B0(a[4]), .B1(n40), .Y(n32) );
  INVX1 U19 ( .A(n29), .Y(N18) );
  AOI22X1 U20 ( .A0(b[1]), .A1(n41), .B0(a[1]), .B1(n40), .Y(n29) );
  INVX1 U21 ( .A(n30), .Y(N19) );
  INVX1 U22 ( .A(n34), .Y(N23) );
  AOI22X1 U23 ( .A0(b[6]), .A1(n41), .B0(a[6]), .B1(n40), .Y(n34) );
  INVX1 U24 ( .A(n35), .Y(N24) );
  INVX1 U25 ( .A(n36), .Y(N25) );
  AOI22X1 U26 ( .A0(b[8]), .A1(n41), .B0(a[8]), .B1(n40), .Y(n36) );
  INVX1 U27 ( .A(n38), .Y(N27) );
  AOI22X1 U28 ( .A0(b[10]), .A1(n41), .B0(a[10]), .B1(n40), .Y(n38) );
  INVX1 U29 ( .A(n42), .Y(N29) );
  AOI22X1 U30 ( .A0(b[12]), .A1(n41), .B0(a[12]), .B1(n40), .Y(n42) );
  AOI22XL U31 ( .A0(b[3]), .A1(n41), .B0(a[3]), .B1(n40), .Y(n31) );
endmodule


module mux13_13_1 ( a, b, sel, enable, out, clk, reset );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel, enable, clk, reset;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N83,
         n3, n6, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42;

  EDFFX4 \out_reg[12]  ( .D(N29), .E(N83), .CK(clk), .Q(out[12]) );
  EDFFX4 \out_reg[11]  ( .D(N28), .E(N83), .CK(clk), .Q(out[11]) );
  EDFFX4 \out_reg[10]  ( .D(N27), .E(N83), .CK(clk), .Q(out[10]) );
  EDFFX4 \out_reg[9]  ( .D(N26), .E(N83), .CK(clk), .Q(out[9]) );
  EDFFX4 \out_reg[8]  ( .D(N25), .E(N83), .CK(clk), .Q(out[8]) );
  EDFFX4 \out_reg[7]  ( .D(N24), .E(N83), .CK(clk), .Q(out[7]) );
  EDFFX4 \out_reg[6]  ( .D(N23), .E(N83), .CK(clk), .Q(out[6]) );
  EDFFX4 \out_reg[5]  ( .D(N22), .E(N83), .CK(clk), .Q(out[5]) );
  EDFFX4 \out_reg[3]  ( .D(N20), .E(N83), .CK(clk), .Q(out[3]) );
  EDFFX4 \out_reg[2]  ( .D(N19), .E(N83), .CK(clk), .Q(out[2]) );
  EDFFX4 \out_reg[0]  ( .D(N17), .E(N83), .CK(clk), .Q(out[0]) );
  DFFHQX4 \out_reg[1]  ( .D(n3), .CK(clk), .Q(out[1]) );
  EDFFX4 \out_reg[4]  ( .D(N21), .E(N83), .CK(clk), .Q(out[4]) );
  INVXL U3 ( .A(n37), .Y(N26) );
  AOI22XL U4 ( .A0(b[1]), .A1(n41), .B0(a[1]), .B1(n40), .Y(n29) );
  AOI22XL U5 ( .A0(b[5]), .A1(n41), .B0(a[5]), .B1(n40), .Y(n33) );
  AOI22XL U6 ( .A0(b[8]), .A1(n41), .B0(a[8]), .B1(n40), .Y(n36) );
  AOI22XL U7 ( .A0(b[10]), .A1(n41), .B0(a[10]), .B1(n40), .Y(n38) );
  AOI22XL U8 ( .A0(b[11]), .A1(n41), .B0(a[11]), .B1(n40), .Y(n39) );
  INVX1 U9 ( .A(n6), .Y(N17) );
  INVX1 U10 ( .A(n42), .Y(N29) );
  INVX1 U11 ( .A(n29), .Y(N18) );
  AOI22XL U12 ( .A0(b[7]), .A1(n41), .B0(a[7]), .B1(n40), .Y(n35) );
  INVX1 U13 ( .A(n34), .Y(N23) );
  INVX1 U14 ( .A(n30), .Y(N19) );
  AOI22X1 U15 ( .A0(b[2]), .A1(n41), .B0(a[2]), .B1(n40), .Y(n30) );
  INVX1 U16 ( .A(n32), .Y(N21) );
  AOI22XL U17 ( .A0(b[4]), .A1(n41), .B0(a[4]), .B1(n40), .Y(n32) );
  INVX1 U18 ( .A(n33), .Y(N22) );
  INVX1 U19 ( .A(n36), .Y(N25) );
  INVX1 U20 ( .A(n38), .Y(N27) );
  NOR2BX1 U21 ( .AN(reset), .B(sel), .Y(n41) );
  AND2X2 U22 ( .A(sel), .B(reset), .Y(n40) );
  NAND2BX1 U23 ( .AN(enable), .B(reset), .Y(N83) );
  INVX1 U24 ( .A(n31), .Y(N20) );
  AOI22X1 U25 ( .A0(b[3]), .A1(n41), .B0(a[3]), .B1(n40), .Y(n31) );
  MX2XL U26 ( .A(out[1]), .B(N18), .S0(N83), .Y(n3) );
  AOI22X1 U27 ( .A0(b[9]), .A1(n41), .B0(a[9]), .B1(n40), .Y(n37) );
  INVX1 U28 ( .A(n39), .Y(N28) );
  AOI22X1 U29 ( .A0(b[6]), .A1(n41), .B0(a[6]), .B1(n40), .Y(n34) );
  INVX1 U30 ( .A(n35), .Y(N24) );
  AOI22XL U31 ( .A0(b[12]), .A1(n41), .B0(a[12]), .B1(n40), .Y(n42) );
  AOI22XL U32 ( .A0(b[0]), .A1(n41), .B0(a[0]), .B1(n40), .Y(n6) );
endmodule


module mux13_13_0 ( a, b, sel, enable, out, clk, reset );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel, enable, clk, reset;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N83,
         n14, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42;

  EDFFX4 \out_reg[1]  ( .D(N18), .E(N83), .CK(clk), .Q(out[1]) );
  EDFFXL \out_reg[10]  ( .D(N27), .E(N83), .CK(clk), .Q(out[10]) );
  EDFFXL \out_reg[8]  ( .D(N25), .E(N83), .CK(clk), .Q(out[8]) );
  EDFFX1 \out_reg[7]  ( .D(N24), .E(N83), .CK(clk), .Q(out[7]) );
  EDFFX1 \out_reg[6]  ( .D(N23), .E(N83), .CK(clk), .Q(out[6]) );
  EDFFX1 \out_reg[4]  ( .D(N21), .E(N83), .CK(clk), .Q(out[4]) );
  EDFFX1 \out_reg[2]  ( .D(N19), .E(N83), .CK(clk), .Q(out[2]) );
  EDFFXL \out_reg[5]  ( .D(N22), .E(N83), .CK(clk), .Q(out[5]) );
  EDFFXL \out_reg[3]  ( .D(N20), .E(N83), .CK(clk), .Q(out[3]) );
  EDFFX1 \out_reg[0]  ( .D(N17), .E(N83), .CK(clk), .Q(out[0]) );
  EDFFX2 \out_reg[12]  ( .D(N29), .E(N83), .CK(clk), .Q(out[12]) );
  EDFFX2 \out_reg[11]  ( .D(N28), .E(N83), .CK(clk), .Q(out[11]) );
  EDFFX2 \out_reg[9]  ( .D(N26), .E(N83), .CK(clk), .Q(out[9]) );
  AOI22XL U3 ( .A0(b[3]), .A1(n41), .B0(a[3]), .B1(n40), .Y(n31) );
  INVXL U4 ( .A(n35), .Y(N24) );
  INVXL U5 ( .A(n34), .Y(N23) );
  AOI22XL U6 ( .A0(b[5]), .A1(n41), .B0(a[5]), .B1(n40), .Y(n33) );
  INVX1 U7 ( .A(n37), .Y(N26) );
  AOI22X1 U8 ( .A0(b[9]), .A1(n41), .B0(a[9]), .B1(n40), .Y(n37) );
  INVX1 U9 ( .A(n39), .Y(N28) );
  AOI22X1 U10 ( .A0(b[11]), .A1(n41), .B0(a[11]), .B1(n40), .Y(n39) );
  INVX1 U11 ( .A(n29), .Y(N18) );
  AOI22X1 U12 ( .A0(b[1]), .A1(n41), .B0(a[1]), .B1(n40), .Y(n29) );
  INVX1 U13 ( .A(n36), .Y(N25) );
  AOI22X1 U14 ( .A0(b[8]), .A1(n41), .B0(a[8]), .B1(n40), .Y(n36) );
  INVX1 U15 ( .A(n38), .Y(N27) );
  AOI22X1 U16 ( .A0(b[10]), .A1(n41), .B0(a[10]), .B1(n40), .Y(n38) );
  INVX1 U17 ( .A(n14), .Y(N17) );
  AOI22X1 U18 ( .A0(b[0]), .A1(n41), .B0(a[0]), .B1(n40), .Y(n14) );
  INVX1 U19 ( .A(n31), .Y(N20) );
  INVX1 U20 ( .A(n32), .Y(N21) );
  AOI22X1 U21 ( .A0(b[4]), .A1(n41), .B0(a[4]), .B1(n40), .Y(n32) );
  INVX1 U22 ( .A(n33), .Y(N22) );
  AOI22X1 U23 ( .A0(b[6]), .A1(n41), .B0(a[6]), .B1(n40), .Y(n34) );
  AOI22X1 U24 ( .A0(b[7]), .A1(n41), .B0(a[7]), .B1(n40), .Y(n35) );
  NAND2BX1 U25 ( .AN(enable), .B(reset), .Y(N83) );
  INVX1 U26 ( .A(n30), .Y(N19) );
  AOI22X1 U27 ( .A0(b[2]), .A1(n41), .B0(a[2]), .B1(n40), .Y(n30) );
  INVX1 U28 ( .A(n42), .Y(N29) );
  AOI22X1 U29 ( .A0(b[12]), .A1(n41), .B0(a[12]), .B1(n40), .Y(n42) );
  NOR2BX1 U30 ( .AN(reset), .B(sel), .Y(n41) );
  AND2X2 U31 ( .A(sel), .B(reset), .Y(n40) );
endmodule


module mux_13_2to1_2 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18;

  INVX1 U1 ( .A(n2), .Y(n3) );
  INVX1 U2 ( .A(n1), .Y(n4) );
  INVX1 U3 ( .A(n2), .Y(n1) );
  INVX1 U4 ( .A(sel), .Y(n2) );
  INVX1 U5 ( .A(n5), .Y(out[0]) );
  AOI22X1 U6 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n2), .Y(n5) );
  INVX1 U7 ( .A(n9), .Y(out[1]) );
  AOI22X1 U8 ( .A0(a[1]), .A1(n3), .B0(b[1]), .B1(n4), .Y(n9) );
  INVX1 U9 ( .A(n10), .Y(out[2]) );
  AOI22X1 U10 ( .A0(a[2]), .A1(n3), .B0(b[2]), .B1(n4), .Y(n10) );
  INVX1 U11 ( .A(n11), .Y(out[3]) );
  AOI22X1 U12 ( .A0(a[3]), .A1(n3), .B0(b[3]), .B1(n4), .Y(n11) );
  INVX1 U13 ( .A(n12), .Y(out[4]) );
  AOI22X1 U14 ( .A0(a[4]), .A1(n3), .B0(b[4]), .B1(n4), .Y(n12) );
  INVX1 U15 ( .A(n13), .Y(out[5]) );
  AOI22X1 U16 ( .A0(a[5]), .A1(n3), .B0(b[5]), .B1(n2), .Y(n13) );
  INVX1 U17 ( .A(n14), .Y(out[6]) );
  AOI22X1 U18 ( .A0(a[6]), .A1(n3), .B0(b[6]), .B1(n4), .Y(n14) );
  INVX1 U19 ( .A(n15), .Y(out[7]) );
  AOI22X1 U20 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n2), .Y(n15) );
  INVX1 U21 ( .A(n17), .Y(out[8]) );
  AOI22X1 U22 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n17) );
  INVX1 U23 ( .A(n18), .Y(out[9]) );
  AOI22X1 U24 ( .A0(n1), .A1(a[9]), .B0(b[9]), .B1(n4), .Y(n18) );
  INVX1 U25 ( .A(n6), .Y(out[10]) );
  AOI22X1 U26 ( .A0(a[10]), .A1(n3), .B0(b[10]), .B1(n2), .Y(n6) );
  INVX1 U27 ( .A(n7), .Y(out[11]) );
  AOI22X1 U28 ( .A0(a[11]), .A1(n3), .B0(b[11]), .B1(n2), .Y(n7) );
  INVX1 U29 ( .A(n8), .Y(out[12]) );
  AOI22X1 U30 ( .A0(a[12]), .A1(n3), .B0(b[12]), .B1(n2), .Y(n8) );
endmodule


module mux_13_2to1_1 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  INVX1 U1 ( .A(n3), .Y(n1) );
  INVX1 U2 ( .A(sel), .Y(n3) );
  INVX1 U3 ( .A(sel), .Y(n2) );
  INVX1 U4 ( .A(n4), .Y(out[0]) );
  AOI22X1 U5 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n4) );
  INVX1 U6 ( .A(n8), .Y(out[1]) );
  AOI22X1 U7 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n2), .Y(n8) );
  INVX1 U8 ( .A(n9), .Y(out[2]) );
  AOI22X1 U9 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n3), .Y(n9) );
  INVX1 U10 ( .A(n10), .Y(out[3]) );
  AOI22X1 U11 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n3), .Y(n10) );
  INVX1 U12 ( .A(n11), .Y(out[4]) );
  AOI22X1 U13 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n2), .Y(n11) );
  INVX1 U14 ( .A(n12), .Y(out[5]) );
  AOI22X1 U15 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n12) );
  INVX1 U16 ( .A(n13), .Y(out[6]) );
  AOI22X1 U17 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n2), .Y(n13) );
  INVX1 U18 ( .A(n14), .Y(out[7]) );
  AOI22X1 U19 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n2), .Y(n14) );
  INVX1 U20 ( .A(n15), .Y(out[8]) );
  AOI22X1 U21 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n2), .Y(n15) );
  INVX1 U22 ( .A(n17), .Y(out[9]) );
  AOI22X1 U23 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n17) );
  INVX1 U24 ( .A(n5), .Y(out[10]) );
  AOI22X1 U25 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n3), .Y(n5) );
  INVX1 U26 ( .A(n6), .Y(out[11]) );
  AOI22X1 U27 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n3), .Y(n6) );
  INVX1 U28 ( .A(n7), .Y(out[12]) );
  AOI22X1 U29 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n2), .Y(n7) );
endmodule


module mux_13_2to1_0 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17
;

  INVX1 U1 ( .A(n3), .Y(n1) );
  INVX1 U2 ( .A(sel), .Y(n3) );
  INVX1 U3 ( .A(sel), .Y(n2) );
  INVX1 U4 ( .A(n4), .Y(out[0]) );
  AOI22X1 U5 ( .A0(a[0]), .A1(n1), .B0(b[0]), .B1(n2), .Y(n4) );
  INVX1 U6 ( .A(n8), .Y(out[1]) );
  AOI22X1 U7 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n3), .Y(n8) );
  INVX1 U8 ( .A(n9), .Y(out[2]) );
  AOI22X1 U9 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n3), .Y(n9) );
  INVX1 U10 ( .A(n10), .Y(out[3]) );
  AOI22X1 U11 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n3), .Y(n10) );
  INVX1 U12 ( .A(n11), .Y(out[4]) );
  AOI22X1 U13 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n2), .Y(n11) );
  INVX1 U14 ( .A(n12), .Y(out[5]) );
  AOI22X1 U15 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n12) );
  INVX1 U16 ( .A(n13), .Y(out[6]) );
  AOI22X1 U17 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n2), .Y(n13) );
  INVX1 U18 ( .A(n14), .Y(out[7]) );
  AOI22X1 U19 ( .A0(a[7]), .A1(sel), .B0(b[7]), .B1(n2), .Y(n14) );
  INVX1 U20 ( .A(n15), .Y(out[8]) );
  AOI22X1 U21 ( .A0(a[8]), .A1(sel), .B0(b[8]), .B1(n2), .Y(n15) );
  INVX1 U22 ( .A(n17), .Y(out[9]) );
  AOI22X1 U23 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n17) );
  INVX1 U24 ( .A(n5), .Y(out[10]) );
  AOI22X1 U25 ( .A0(a[10]), .A1(n1), .B0(b[10]), .B1(n2), .Y(n5) );
  INVX1 U26 ( .A(n6), .Y(out[11]) );
  AOI22X1 U27 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n2), .Y(n6) );
  INVX1 U28 ( .A(n7), .Y(out[12]) );
  AOI22X1 U29 ( .A0(a[12]), .A1(n1), .B0(b[12]), .B1(n3), .Y(n7) );
endmodule


module multiplier_14 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n36, n37, n38, n39, n43, n47, n49, n50, n51, n52,
         n53, n54, n55, n57, n58, n59, n61, n63, n64, n77, n81, n83, n84, n85,
         n86, n87, n92, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n122, n127, n128, n131,
         n132, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n202, n203, n204, n205, n210, n211,
         n212, n213, n214, n215, n216, n217, n219, n220, n221, n239, n240,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n259, n260,
         n261, n262, n263, n264, n265, n266, n286, n288, n289, n290, n291,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n311, n314, n315, n316, n317, n318, n319, n320, n321, n323, n324,
         n325, n326, n327, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527;

  OAI21X1 U1 ( .A0(n368), .A1(n367), .B0(n366), .Y(n436) );
  NOR2X1 U2 ( .A(n365), .B(n23), .Y(n211) );
  NOR2X1 U3 ( .A(n365), .B(n22), .Y(n290) );
  OAI21XL U4 ( .A0(n85), .A1(n29), .B0(n360), .Y(n213) );
  OAI211X1 U5 ( .A0(n178), .A1(n29), .B0(n28), .C0(n81), .Y(n165) );
  OAI221XL U6 ( .A0(n29), .A1(n53), .B0(n52), .B1(n365), .C0(n361), .Y(n362)
         );
  NOR2X1 U7 ( .A(n365), .B(n377), .Y(n57) );
  XNOR3X2 U8 ( .A(n370), .B(n453), .C(n175), .Y(c[2]) );
  NOR2X1 U9 ( .A(n29), .B(n22), .Y(n303) );
  NOR2X1 U10 ( .A(n508), .B(n10), .Y(n399) );
  XOR3X2 U11 ( .A(n338), .B(n326), .C(n337), .Y(c[10]) );
  NAND2BX1 U12 ( .AN(a[12]), .B(a[11]), .Y(n163) );
  INVX1 U13 ( .A(a[12]), .Y(n365) );
  BUFX4 U14 ( .A(b[4]), .Y(n81) );
  CLKINVX3 U15 ( .A(n138), .Y(n321) );
  NOR2X1 U16 ( .A(n363), .B(n380), .Y(n364) );
  XOR2X1 U17 ( .A(n452), .B(n451), .Y(n481) );
  INVX1 U18 ( .A(n373), .Y(n369) );
  XOR2X1 U19 ( .A(n104), .B(n64), .Y(n138) );
  AOI21X1 U20 ( .A0(n25), .A1(n103), .B0(n102), .Y(n104) );
  INVX1 U21 ( .A(n481), .Y(n372) );
  NAND2BX2 U22 ( .AN(a[12]), .B(a[11]), .Y(n360) );
  NAND2X1 U23 ( .A(n9), .B(n27), .Y(n51) );
  INVX2 U24 ( .A(b[10]), .Y(n26) );
  OAI2BB1XL U25 ( .A0N(a[11]), .A1N(n81), .B0(n380), .Y(n366) );
  INVX1 U26 ( .A(b[3]), .Y(n380) );
  XNOR3X2 U27 ( .A(n371), .B(n478), .C(n370), .Y(n47) );
  XOR2X1 U28 ( .A(n527), .B(n50), .Y(n346) );
  INVX1 U29 ( .A(n365), .Y(n28) );
  INVX1 U30 ( .A(n302), .Y(n367) );
  INVX1 U31 ( .A(a[11]), .Y(n29) );
  BUFX3 U32 ( .A(b[3]), .Y(n1) );
  BUFX3 U33 ( .A(n53), .Y(n2) );
  NAND2X1 U34 ( .A(b[1]), .B(n521), .Y(n53) );
  NAND2X1 U35 ( .A(b[0]), .B(n520), .Y(n3) );
  NAND2X1 U36 ( .A(b[0]), .B(n520), .Y(n52) );
  INVX1 U37 ( .A(b[0]), .Y(n4) );
  INVX1 U38 ( .A(n378), .Y(n5) );
  INVX1 U39 ( .A(n374), .Y(n6) );
  INVX1 U40 ( .A(n377), .Y(n7) );
  INVX1 U41 ( .A(a[10]), .Y(n8) );
  INVX1 U42 ( .A(n8), .Y(n9) );
  INVX1 U43 ( .A(a[9]), .Y(n10) );
  INVX1 U44 ( .A(n10), .Y(n11) );
  INVX1 U45 ( .A(n10), .Y(n12) );
  INVX1 U46 ( .A(a[8]), .Y(n13) );
  INVX1 U47 ( .A(n13), .Y(n14) );
  INVX1 U48 ( .A(n13), .Y(n15) );
  INVX1 U49 ( .A(a[7]), .Y(n16) );
  INVXL U50 ( .A(n16), .Y(n17) );
  INVX1 U51 ( .A(n507), .Y(n18) );
  INVX1 U52 ( .A(n487), .Y(n19) );
  INVX1 U53 ( .A(n450), .Y(n20) );
  NAND2X1 U54 ( .A(n97), .B(b[11]), .Y(n146) );
  INVX1 U55 ( .A(n519), .Y(n21) );
  BUFX3 U56 ( .A(b[9]), .Y(n22) );
  BUFX3 U57 ( .A(b[8]), .Y(n23) );
  INVX1 U58 ( .A(n246), .Y(n24) );
  AOI21X1 U59 ( .A0(n84), .A1(n181), .B0(n180), .Y(n194) );
  BUFX3 U60 ( .A(b[6]), .Y(n84) );
  XOR2X2 U61 ( .A(n137), .B(n136), .Y(n173) );
  XNOR2XL U62 ( .A(n33), .B(n369), .Y(n262) );
  XOR2X2 U63 ( .A(n34), .B(n170), .Y(n33) );
  OAI21XL U64 ( .A0(n9), .A1(n359), .B0(n53), .Y(n388) );
  OAI21XL U65 ( .A0(n100), .A1(n359), .B0(n53), .Y(n486) );
  NOR2X2 U66 ( .A(n250), .B(n249), .Y(n259) );
  XOR2X4 U67 ( .A(n151), .B(n150), .Y(n370) );
  BUFX3 U68 ( .A(b[11]), .Y(n25) );
  NAND2XL U69 ( .A(n98), .B(n25), .Y(n444) );
  INVXL U70 ( .A(n26), .Y(n27) );
  NAND2XL U71 ( .A(n92), .B(n27), .Y(n332) );
  NAND2XL U72 ( .A(n99), .B(n27), .Y(n445) );
  NAND2XL U73 ( .A(n98), .B(n27), .Y(n429) );
  NAND2XL U74 ( .A(b[10]), .B(n97), .Y(n109) );
  NAND2BXL U75 ( .AN(n85), .B(n28), .Y(n247) );
  NOR2BXL U76 ( .AN(a[12]), .B(n77), .Y(n127) );
  NAND2BX2 U77 ( .AN(a[11]), .B(a[12]), .Y(n302) );
  INVXL U78 ( .A(n29), .Y(n30) );
  INVXL U79 ( .A(n262), .Y(n205) );
  XOR2X1 U80 ( .A(n55), .B(n431), .Y(c[1]) );
  XNOR3X2 U81 ( .A(n55), .B(n205), .C(n204), .Y(c[4]) );
  XOR2X1 U82 ( .A(n480), .B(n479), .Y(c[5]) );
  AOI22XL U83 ( .A0(n17), .A1(n506), .B0(n15), .B1(n505), .Y(n510) );
  AOI2BB2XL U84 ( .B0(b[0]), .B1(n367), .A0N(n360), .A1N(n359), .Y(n361) );
  XNOR2X1 U85 ( .A(n266), .B(n31), .Y(n54) );
  NAND2XL U86 ( .A(n99), .B(n25), .Y(n457) );
  NAND2XL U87 ( .A(n97), .B(n1), .Y(n491) );
  NAND2XL U88 ( .A(n98), .B(n1), .Y(n500) );
  NAND2XL U89 ( .A(n14), .B(n83), .Y(n58) );
  NAND2XL U90 ( .A(n1), .B(n18), .Y(n526) );
  INVXL U91 ( .A(n358), .Y(n174) );
  XOR3X2 U92 ( .A(n32), .B(n259), .C(n254), .Y(n31) );
  XNOR2X1 U93 ( .A(n240), .B(n239), .Y(n32) );
  XOR3X2 U94 ( .A(n454), .B(n455), .C(n152), .Y(n34) );
  NOR2XL U95 ( .A(n374), .B(n378), .Y(n403) );
  NOR2XL U96 ( .A(n376), .B(n380), .Y(n458) );
  NOR2XL U97 ( .A(n375), .B(n378), .Y(n501) );
  XNOR2X1 U98 ( .A(n481), .B(n371), .Y(n175) );
  XOR3X2 U99 ( .A(n36), .B(n390), .C(n37), .Y(n337) );
  XOR3X2 U100 ( .A(n391), .B(n330), .C(n327), .Y(n36) );
  XNOR3X2 U101 ( .A(n336), .B(n335), .C(n334), .Y(n37) );
  XNOR2X1 U102 ( .A(n321), .B(n57), .Y(n358) );
  AOI22XL U103 ( .A0(n87), .A1(n106), .B0(n25), .B1(n105), .Y(n371) );
  NAND2XL U104 ( .A(n85), .B(n100), .Y(n383) );
  AOI21XL U105 ( .A0(n30), .A1(n164), .B0(n363), .Y(n166) );
  NAND2XL U106 ( .A(n22), .B(n9), .Y(n215) );
  NAND2XL U107 ( .A(n5), .B(n97), .Y(n330) );
  NAND2XL U108 ( .A(a[7]), .B(n22), .Y(n455) );
  NAND2XL U109 ( .A(n85), .B(n15), .Y(n438) );
  AOI22XL U110 ( .A0(n15), .A1(n523), .B0(n12), .B1(n522), .Y(n524) );
  NAND2XL U111 ( .A(n14), .B(n87), .Y(n288) );
  NAND2XL U112 ( .A(n11), .B(b[11]), .Y(n286) );
  NAND2XL U113 ( .A(b[8]), .B(n14), .Y(n162) );
  NAND2XL U114 ( .A(n85), .B(n11), .Y(n153) );
  NAND2XL U115 ( .A(n98), .B(n86), .Y(n385) );
  NAND2XL U116 ( .A(n99), .B(b[8]), .Y(n386) );
  NAND2XL U117 ( .A(n87), .B(n96), .Y(n147) );
  OAI21XL U118 ( .A0(n303), .A1(n363), .B0(n27), .Y(n304) );
  NAND2BXL U119 ( .AN(n84), .B(n28), .Y(n179) );
  INVXL U120 ( .A(n85), .Y(n378) );
  NAND2XL U121 ( .A(n17), .B(n7), .Y(n219) );
  NAND2XL U122 ( .A(n15), .B(n27), .Y(n251) );
  XNOR3X2 U123 ( .A(n38), .B(n396), .C(n306), .Y(n527) );
  NAND2XL U124 ( .A(n12), .B(n87), .Y(n38) );
  OAI2BB1X1 U125 ( .A0N(a[11]), .A1N(n26), .B0(n360), .Y(n103) );
  OAI2BB1X1 U126 ( .A0N(b[3]), .A1N(n142), .B0(n141), .Y(n144) );
  NAND2XL U127 ( .A(n360), .B(n139), .Y(n142) );
  NAND2XL U128 ( .A(b[4]), .B(n17), .Y(n401) );
  NAND2XL U129 ( .A(n97), .B(b[4]), .Y(n499) );
  NAND2XL U130 ( .A(n81), .B(n99), .Y(n525) );
  XNOR3X2 U131 ( .A(n323), .B(n321), .C(n524), .Y(n324) );
  NAND2XL U132 ( .A(n92), .B(n22), .Y(n319) );
  NAND2XL U133 ( .A(n85), .B(n96), .Y(n318) );
  NAND2XL U134 ( .A(n77), .B(n9), .Y(n407) );
  NAND2XL U135 ( .A(n9), .B(n1), .Y(n135) );
  NAND2XL U136 ( .A(n100), .B(n27), .Y(n454) );
  NAND2XL U137 ( .A(n84), .B(n18), .Y(n404) );
  NAND2XL U138 ( .A(n97), .B(n83), .Y(n503) );
  NAND2XL U139 ( .A(n24), .B(n96), .Y(n502) );
  NAND2XL U140 ( .A(n81), .B(n15), .Y(n408) );
  NAND2XL U141 ( .A(n98), .B(b[4]), .Y(n511) );
  NAND2XL U142 ( .A(n100), .B(n86), .Y(n442) );
  NAND2XL U143 ( .A(n20), .B(n23), .Y(n395) );
  NAND2XL U144 ( .A(n23), .B(n95), .Y(n311) );
  NAND2XL U145 ( .A(n100), .B(n25), .Y(n468) );
  NAND2XL U146 ( .A(n92), .B(n5), .Y(n264) );
  NAND2XL U147 ( .A(n24), .B(n92), .Y(n482) );
  NAND2XL U148 ( .A(n15), .B(n25), .Y(n217) );
  XOR2X1 U149 ( .A(n191), .B(n190), .Y(n192) );
  NAND2XL U150 ( .A(a[10]), .B(n87), .Y(n64) );
  NAND2XL U151 ( .A(n83), .B(n9), .Y(n437) );
  NAND2XL U152 ( .A(n99), .B(n87), .Y(n189) );
  NAND2XL U153 ( .A(n86), .B(n14), .Y(n188) );
  NAND2XL U154 ( .A(n98), .B(n87), .Y(n456) );
  NAND2XL U155 ( .A(n84), .B(n97), .Y(n314) );
  NAND2XL U156 ( .A(n21), .B(n22), .Y(n394) );
  NAND2XL U157 ( .A(b[5]), .B(n95), .Y(n483) );
  NAND2XL U158 ( .A(a[7]), .B(n27), .Y(n469) );
  NAND2XL U159 ( .A(n98), .B(n24), .Y(n331) );
  NAND2XL U160 ( .A(n22), .B(n95), .Y(n333) );
  NAND2XL U161 ( .A(n84), .B(n17), .Y(n384) );
  NAND2XL U162 ( .A(n85), .B(a[7]), .Y(n428) );
  NAND2XL U163 ( .A(n1), .B(n17), .Y(n393) );
  NAND2XL U164 ( .A(n81), .B(n100), .Y(n392) );
  NAND2XL U165 ( .A(n6), .B(n83), .Y(n327) );
  NAND2BXL U166 ( .AN(b[11]), .B(a[12]), .Y(n101) );
  NAND2XL U167 ( .A(n1), .B(n12), .Y(n409) );
  NAND2XL U168 ( .A(a[7]), .B(n23), .Y(n443) );
  NAND2XL U169 ( .A(n96), .B(n81), .Y(n490) );
  NAND2XL U170 ( .A(n85), .B(a[10]), .Y(n187) );
  NAND2XL U171 ( .A(b[8]), .B(n11), .Y(n182) );
  AOI22XL U172 ( .A0(n9), .A1(n398), .B0(n30), .B1(n397), .Y(n400) );
  NAND2XL U173 ( .A(n1), .B(n15), .Y(n402) );
  XNOR2X1 U174 ( .A(n39), .B(n315), .Y(n316) );
  NAND2XL U175 ( .A(n17), .B(n77), .Y(n39) );
  XOR3X2 U176 ( .A(n47), .B(n43), .C(n372), .Y(n479) );
  XNOR2XL U177 ( .A(n369), .B(n31), .Y(n43) );
  XOR3X2 U178 ( .A(n49), .B(n299), .C(n326), .Y(n300) );
  NAND2XL U179 ( .A(n24), .B(n95), .Y(n49) );
  NAND2BXL U180 ( .AN(n84), .B(a[11]), .Y(n248) );
  AOI22XL U181 ( .A0(n18), .A1(n496), .B0(n17), .B1(n495), .Y(n498) );
  NAND2XL U182 ( .A(n92), .B(b[4]), .Y(n203) );
  NAND2XL U183 ( .A(n7), .B(n95), .Y(n107) );
  NAND2XL U184 ( .A(b[11]), .B(n96), .Y(n108) );
  NAND2XL U185 ( .A(n84), .B(n14), .Y(n61) );
  NAND2XL U186 ( .A(n11), .B(n83), .Y(n63) );
  NAND2XL U187 ( .A(n12), .B(n81), .Y(n59) );
  INVXL U188 ( .A(n100), .Y(n507) );
  NAND2XL U189 ( .A(n83), .B(n17), .Y(n405) );
  NAND2XL U190 ( .A(n92), .B(n7), .Y(n414) );
  NAND2XL U191 ( .A(n25), .B(n9), .Y(n396) );
  NAND2BXL U192 ( .AN(n77), .B(a[11]), .Y(n139) );
  NAND2XL U193 ( .A(n99), .B(n86), .Y(n430) );
  NAND2XL U194 ( .A(n100), .B(n23), .Y(n427) );
  INVXL U195 ( .A(n87), .Y(n377) );
  INVXL U196 ( .A(n81), .Y(n164) );
  AND2X1 U197 ( .A(a[10]), .B(n81), .Y(n145) );
  AND2X1 U198 ( .A(n84), .B(a[10]), .Y(n169) );
  AND2X1 U199 ( .A(n12), .B(b[10]), .Y(n216) );
  INVX1 U200 ( .A(n163), .Y(n363) );
  AND2X1 U201 ( .A(n98), .B(n83), .Y(n315) );
  XOR3X2 U202 ( .A(n51), .B(n298), .C(n297), .Y(n50) );
  NAND2XL U203 ( .A(n360), .B(n289), .Y(n296) );
  NAND2BXL U204 ( .AN(b[8]), .B(n30), .Y(n289) );
  XOR2X1 U205 ( .A(n441), .B(n440), .Y(n449) );
  XOR2X1 U206 ( .A(n439), .B(n438), .Y(n440) );
  NAND2XL U207 ( .A(n84), .B(n12), .Y(n439) );
  NAND2XL U208 ( .A(n23), .B(n96), .Y(n335) );
  NAND2XL U209 ( .A(n92), .B(n25), .Y(n351) );
  NAND2XL U210 ( .A(n18), .B(b[5]), .Y(n347) );
  NAND2XL U211 ( .A(n6), .B(n24), .Y(n348) );
  NAND2XL U212 ( .A(n19), .B(n5), .Y(n349) );
  NAND2XL U213 ( .A(n20), .B(n22), .Y(n417) );
  NAND2XL U214 ( .A(b[4]), .B(n95), .Y(n474) );
  NAND2XL U215 ( .A(a[1]), .B(n25), .Y(n419) );
  AND2X1 U216 ( .A(n15), .B(n77), .Y(n390) );
  AND2X1 U217 ( .A(n23), .B(a[0]), .Y(n517) );
  NAND2XL U218 ( .A(n1), .B(a[1]), .Y(n195) );
  NAND2XL U219 ( .A(n21), .B(n27), .Y(n420) );
  NAND2XL U220 ( .A(n95), .B(n27), .Y(n350) );
  NAND2XL U221 ( .A(n19), .B(n23), .Y(n418) );
  OAI2BB1X1 U222 ( .A0N(n77), .A1N(n131), .B0(n128), .Y(n134) );
  NAND2XL U223 ( .A(n360), .B(n122), .Y(n131) );
  NAND2BXL U224 ( .AN(b[1]), .B(n30), .Y(n122) );
  INVXL U225 ( .A(b[1]), .Y(n359) );
  XOR2X1 U226 ( .A(n54), .B(n372), .Y(n260) );
  XOR3X2 U227 ( .A(n253), .B(n252), .C(n251), .Y(n254) );
  XOR3X2 U228 ( .A(n346), .B(n517), .C(n518), .Y(c[8]) );
  XNOR3X2 U229 ( .A(n174), .B(n33), .C(n173), .Y(n176) );
  XOR2X1 U230 ( .A(n266), .B(n50), .Y(n326) );
  XOR3X2 U231 ( .A(n501), .B(n31), .C(n373), .Y(n381) );
  XNOR3X2 U232 ( .A(n33), .B(n494), .C(n210), .Y(n261) );
  XOR2X1 U233 ( .A(n484), .B(n57), .Y(n210) );
  XOR2X1 U234 ( .A(n493), .B(n492), .Y(n494) );
  XOR2X1 U235 ( .A(n483), .B(n482), .Y(n484) );
  XOR3X2 U236 ( .A(n354), .B(n353), .C(n352), .Y(n355) );
  XOR2X1 U237 ( .A(n394), .B(n395), .Y(n353) );
  XNOR3X2 U238 ( .A(n401), .B(n351), .C(n350), .Y(n352) );
  XOR2X1 U239 ( .A(n371), .B(n57), .Y(n354) );
  XNOR3X2 U240 ( .A(n169), .B(n168), .C(n167), .Y(n170) );
  XOR2X1 U241 ( .A(n261), .B(n260), .Y(c[6]) );
  XOR2X1 U242 ( .A(n424), .B(n423), .Y(c[12]) );
  XOR2X1 U243 ( .A(n516), .B(n515), .Y(n518) );
  XOR2X1 U244 ( .A(n514), .B(n513), .Y(n515) );
  XOR2X1 U245 ( .A(n381), .B(n504), .Y(n516) );
  XOR2X1 U246 ( .A(n512), .B(n511), .Y(n513) );
  XOR2X1 U247 ( .A(n463), .B(n458), .Y(n177) );
  XOR2X1 U248 ( .A(n462), .B(n461), .Y(n463) );
  NOR2X1 U249 ( .A(n375), .B(n508), .Y(n461) );
  XOR3X2 U250 ( .A(n174), .B(n173), .C(n370), .Y(n55) );
  XNOR2X1 U251 ( .A(n301), .B(n300), .Y(c[7]) );
  XOR3X2 U252 ( .A(n177), .B(n176), .C(n175), .Y(c[3]) );
  XNOR3X2 U253 ( .A(n325), .B(n54), .C(n324), .Y(c[9]) );
  XNOR3X2 U254 ( .A(n357), .B(n356), .C(n355), .Y(c[11]) );
  NOR2X1 U255 ( .A(n508), .B(n374), .Y(n497) );
  OAI21XL U256 ( .A0(n25), .A1(n29), .B0(n360), .Y(n106) );
  OAI21XL U257 ( .A0(n12), .A1(n520), .B0(n2), .Y(n523) );
  OAI21XL U258 ( .A0(n15), .A1(n4), .B0(n52), .Y(n522) );
  MXI2X1 U259 ( .A(n365), .B(n364), .S0(n81), .Y(n368) );
  AOI22X1 U260 ( .A0(n96), .A1(n460), .B0(n97), .B1(n459), .Y(n462) );
  OAI21XL U261 ( .A0(n97), .A1(n359), .B0(n53), .Y(n460) );
  OAI21XL U262 ( .A0(n96), .A1(n4), .B0(n3), .Y(n459) );
  AOI22X1 U263 ( .A0(n9), .A1(n389), .B0(n12), .B1(n388), .Y(n391) );
  OAI21XL U264 ( .A0(n12), .A1(n4), .B0(n3), .Y(n389) );
  AOI21X1 U265 ( .A0(n360), .A1(n248), .B0(n378), .Y(n249) );
  INVXL U266 ( .A(n84), .Y(n246) );
  OAI2BB1X1 U267 ( .A0N(n22), .A1N(n305), .B0(n304), .Y(n306) );
  OAI21XL U268 ( .A0(n15), .A1(n359), .B0(n53), .Y(n506) );
  OAI21XL U269 ( .A0(n19), .A1(n359), .B0(n2), .Y(n465) );
  OAI21XL U270 ( .A0(n17), .A1(n359), .B0(n2), .Y(n496) );
  OAI21XL U271 ( .A0(n30), .A1(n359), .B0(n2), .Y(n398) );
  OAI21XL U272 ( .A0(n99), .A1(n4), .B0(n52), .Y(n485) );
  OAI21XL U273 ( .A0(n17), .A1(n4), .B0(n3), .Y(n505) );
  OAI21XL U274 ( .A0(n95), .A1(n521), .B0(n3), .Y(n432) );
  OAI21XL U275 ( .A0(n20), .A1(n521), .B0(n52), .Y(n464) );
  AOI22X1 U276 ( .A0(n19), .A1(n471), .B0(n6), .B1(n470), .Y(n472) );
  OAI21XL U277 ( .A0(n6), .A1(n359), .B0(n2), .Y(n471) );
  OAI21XL U278 ( .A0(n98), .A1(n4), .B0(n3), .Y(n470) );
  OAI21XL U279 ( .A0(n18), .A1(n4), .B0(n52), .Y(n495) );
  OAI21XL U280 ( .A0(n9), .A1(n4), .B0(n52), .Y(n397) );
  INVX1 U281 ( .A(n77), .Y(n508) );
  OAI21XL U282 ( .A0(n166), .A1(n178), .B0(n165), .Y(n167) );
  XNOR3X2 U283 ( .A(n429), .B(n149), .C(n148), .Y(n150) );
  XNOR3X2 U284 ( .A(n145), .B(n144), .C(n143), .Y(n151) );
  OAI21XL U285 ( .A0(n290), .A1(n367), .B0(n23), .Y(n291) );
  XNOR3X2 U286 ( .A(n383), .B(n111), .C(n110), .Y(n137) );
  XNOR3X2 U287 ( .A(n135), .B(n134), .C(n132), .Y(n136) );
  XNOR3X2 U288 ( .A(n194), .B(n193), .C(n192), .Y(n373) );
  XNOR2X1 U289 ( .A(n469), .B(n468), .Y(n193) );
  XOR2X1 U290 ( .A(n221), .B(n220), .Y(n266) );
  XOR2X1 U291 ( .A(n219), .B(n217), .Y(n220) );
  XNOR3X2 U292 ( .A(n216), .B(n215), .C(n214), .Y(n221) );
  NOR2X1 U293 ( .A(n377), .B(n450), .Y(n451) );
  XOR2X1 U294 ( .A(n449), .B(n448), .Y(n452) );
  INVX1 U295 ( .A(n97), .Y(n450) );
  NAND2X1 U296 ( .A(n100), .B(n87), .Y(n252) );
  NAND2X1 U297 ( .A(a[7]), .B(b[11]), .Y(n239) );
  XOR2X1 U298 ( .A(n491), .B(n490), .Y(n492) );
  XNOR2X1 U299 ( .A(n187), .B(n182), .Y(n191) );
  AND2X2 U300 ( .A(n83), .B(n92), .Y(n478) );
  XOR2X1 U301 ( .A(n265), .B(n264), .Y(n299) );
  NAND2X1 U302 ( .A(b[5]), .B(n96), .Y(n265) );
  OAI2BB1X1 U303 ( .A0N(n22), .A1N(n296), .B0(n291), .Y(n297) );
  XOR2X1 U304 ( .A(n435), .B(n434), .Y(n453) );
  NOR2X1 U305 ( .A(n376), .B(n508), .Y(n434) );
  AOI22X1 U306 ( .A0(n95), .A1(n433), .B0(n21), .B1(n432), .Y(n435) );
  OAI21XL U307 ( .A0(n21), .A1(n359), .B0(n2), .Y(n433) );
  XOR2X1 U308 ( .A(n288), .B(n286), .Y(n298) );
  XOR2X1 U309 ( .A(n162), .B(n153), .Y(n168) );
  XOR2X1 U310 ( .A(n385), .B(n386), .Y(n111) );
  XOR2X1 U311 ( .A(n147), .B(n146), .Y(n149) );
  XOR2X1 U312 ( .A(n189), .B(n188), .Y(n190) );
  XOR2X1 U313 ( .A(n447), .B(n446), .Y(n448) );
  XOR2X1 U314 ( .A(n443), .B(n442), .Y(n447) );
  XOR2X1 U315 ( .A(n445), .B(n444), .Y(n446) );
  XOR2X1 U316 ( .A(n411), .B(n410), .Y(n412) );
  XOR2X1 U317 ( .A(n409), .B(n408), .Y(n410) );
  XOR2X1 U318 ( .A(n362), .B(n407), .Y(n411) );
  XNOR3X2 U319 ( .A(n498), .B(n263), .C(n262), .Y(n301) );
  XOR3X2 U320 ( .A(n499), .B(n500), .C(n497), .Y(n263) );
  OAI2BB1X1 U321 ( .A0N(n30), .A1N(n178), .B0(n360), .Y(n181) );
  XNOR3X2 U322 ( .A(n400), .B(n346), .C(n339), .Y(n357) );
  XNOR2X1 U323 ( .A(n399), .B(n402), .Y(n339) );
  NAND2X1 U324 ( .A(a[10]), .B(b[8]), .Y(n240) );
  XNOR3X2 U325 ( .A(n317), .B(n316), .C(n527), .Y(n325) );
  XOR2X1 U326 ( .A(n314), .B(n311), .Y(n317) );
  XNOR3X2 U327 ( .A(n58), .B(n59), .C(n384), .Y(n132) );
  XNOR3X2 U328 ( .A(n61), .B(n63), .C(n428), .Y(n143) );
  XOR3X2 U329 ( .A(n525), .B(n526), .C(n320), .Y(n323) );
  XNOR3X2 U330 ( .A(n467), .B(n203), .C(n202), .Y(n204) );
  XOR2X1 U331 ( .A(n195), .B(n466), .Y(n202) );
  AOI22X1 U332 ( .A0(n20), .A1(n465), .B0(n19), .B1(n464), .Y(n467) );
  XNOR3X2 U333 ( .A(n109), .B(n108), .C(n107), .Y(n110) );
  NAND2X1 U334 ( .A(n86), .B(n11), .Y(n253) );
  XNOR3X2 U335 ( .A(n387), .B(n338), .C(n173), .Y(c[0]) );
  XOR2X1 U336 ( .A(n489), .B(n488), .Y(n493) );
  NOR2X1 U337 ( .A(n508), .B(n487), .Y(n488) );
  AOI22X1 U338 ( .A0(n99), .A1(n486), .B0(n100), .B1(n485), .Y(n489) );
  INVX1 U339 ( .A(n98), .Y(n487) );
  XOR2X1 U340 ( .A(n510), .B(n509), .Y(n514) );
  NOR2X1 U341 ( .A(n508), .B(n507), .Y(n509) );
  XOR2X1 U342 ( .A(n416), .B(n415), .Y(n424) );
  XNOR2X1 U343 ( .A(n414), .B(n527), .Y(n415) );
  XOR2X1 U344 ( .A(n413), .B(n412), .Y(n416) );
  XOR2X1 U345 ( .A(n436), .B(n437), .Y(n441) );
  XOR2X1 U346 ( .A(n382), .B(n406), .Y(n413) );
  XOR2X1 U347 ( .A(n405), .B(n404), .Y(n406) );
  XOR2X1 U348 ( .A(n358), .B(n403), .Y(n382) );
  XOR2X1 U349 ( .A(n477), .B(n476), .Y(n480) );
  XOR2X1 U350 ( .A(n475), .B(n474), .Y(n476) );
  XOR2X1 U351 ( .A(n473), .B(n472), .Y(n477) );
  NAND2X1 U352 ( .A(n21), .B(n1), .Y(n475) );
  INVX1 U353 ( .A(n99), .Y(n374) );
  OAI2BB1X1 U354 ( .A0N(n23), .A1N(n213), .B0(n212), .Y(n214) );
  OAI21XL U355 ( .A0(n211), .A1(n367), .B0(n85), .Y(n212) );
  OAI21XL U356 ( .A0(n140), .A1(n367), .B0(n77), .Y(n141) );
  NOR2BX1 U357 ( .AN(a[12]), .B(b[3]), .Y(n140) );
  XNOR2X1 U358 ( .A(n430), .B(n427), .Y(n148) );
  INVX1 U359 ( .A(n83), .Y(n178) );
  XOR2X1 U360 ( .A(n456), .B(n457), .Y(n152) );
  AOI22X1 U361 ( .A0(a[0]), .A1(n426), .B0(a[1]), .B1(n425), .Y(n431) );
  OAI21XL U362 ( .A0(a[1]), .A1(n520), .B0(n2), .Y(n426) );
  OAI21XL U363 ( .A0(n92), .A1(n4), .B0(n3), .Y(n425) );
  NOR2X1 U364 ( .A(n508), .B(n519), .Y(n466) );
  INVX1 U365 ( .A(n96), .Y(n519) );
  NOR2X1 U366 ( .A(n376), .B(n4), .Y(n387) );
  XOR2X1 U367 ( .A(n503), .B(n502), .Y(n504) );
  XOR2X1 U368 ( .A(n422), .B(n421), .Y(n423) );
  XOR2X1 U369 ( .A(n418), .B(n417), .Y(n422) );
  XOR2X1 U370 ( .A(n420), .B(n419), .Y(n421) );
  NAND2X1 U371 ( .A(n99), .B(n1), .Y(n512) );
  NAND2X1 U372 ( .A(n20), .B(n77), .Y(n473) );
  XOR3X2 U373 ( .A(n333), .B(n332), .C(n331), .Y(n334) );
  XNOR3X2 U374 ( .A(n349), .B(n348), .C(n347), .Y(n356) );
  INVX1 U375 ( .A(n92), .Y(n376) );
  XOR2X1 U376 ( .A(n319), .B(n318), .Y(n320) );
  XOR2X1 U377 ( .A(n393), .B(n392), .Y(n336) );
  INVX1 U378 ( .A(n95), .Y(n375) );
  BUFX3 U379 ( .A(a[3]), .Y(n97) );
  BUFX3 U380 ( .A(a[6]), .Y(n100) );
  BUFX3 U381 ( .A(a[2]), .Y(n96) );
  BUFX3 U382 ( .A(a[4]), .Y(n98) );
  BUFX3 U383 ( .A(a[5]), .Y(n99) );
  BUFX3 U384 ( .A(b[9]), .Y(n86) );
  BUFX3 U385 ( .A(a[1]), .Y(n95) );
  BUFX3 U386 ( .A(b[12]), .Y(n87) );
  BUFX3 U387 ( .A(b[7]), .Y(n85) );
  INVX1 U388 ( .A(b[0]), .Y(n521) );
  INVX1 U389 ( .A(b[1]), .Y(n520) );
  BUFX3 U390 ( .A(b[5]), .Y(n83) );
  BUFX3 U391 ( .A(b[2]), .Y(n77) );
  OAI21XL U392 ( .A0(n127), .A1(n367), .B0(b[1]), .Y(n128) );
  BUFX3 U393 ( .A(a[0]), .Y(n92) );
  OAI21XL U394 ( .A0(n87), .A1(n365), .B0(n302), .Y(n105) );
  OAI2BB1X1 U395 ( .A0N(n28), .A1N(n26), .B0(n302), .Y(n305) );
  AOI21X1 U396 ( .A0(n302), .A1(n179), .B0(n178), .Y(n180) );
  AOI21X1 U397 ( .A0(n302), .A1(n247), .B0(n246), .Y(n250) );
  AOI21X1 U398 ( .A0(n302), .A1(n101), .B0(n26), .Y(n102) );
  XOR2X1 U399 ( .A(n138), .B(n371), .Y(n338) );
endmodule


module multiplier_13 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n47, n49, n50, n51, n52,
         n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n92, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n122, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n202, n203,
         n204, n205, n210, n211, n212, n213, n214, n215, n216, n217, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n230, n233,
         n234, n235, n236, n237, n238, n239, n240, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n259, n260, n261, n262, n263, n264,
         n265, n266, n278, n280, n286, n288, n289, n290, n291, n292, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n343, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507;

  XOR2X2 U1 ( .A(n291), .B(n180), .Y(n215) );
  AOI22XL U2 ( .A0(n25), .A1(n467), .B0(a[5]), .B1(n466), .Y(n468) );
  AND2X1 U3 ( .A(a[10]), .B(n13), .Y(n128) );
  XOR2X1 U4 ( .A(n167), .B(n166), .Y(n181) );
  NAND3X1 U5 ( .A(n335), .B(n334), .C(n333), .Y(n394) );
  OAI21XL U6 ( .A0(n1), .A1(n102), .B0(n325), .Y(n326) );
  INVX1 U7 ( .A(n111), .Y(n1) );
  OAI21XL U8 ( .A0(n386), .A1(n122), .B0(n102), .Y(n126) );
  AOI21X1 U9 ( .A0(n37), .A1(n110), .B0(n2), .Y(n64) );
  INVX1 U10 ( .A(n385), .Y(n2) );
  OAI2BB1X1 U11 ( .A0N(n103), .A1N(n127), .B0(n126), .Y(n129) );
  OAI211X1 U12 ( .A0(n3), .A1(n65), .B0(n388), .C0(n387), .Y(n389) );
  INVX1 U13 ( .A(n35), .Y(n3) );
  OAI21XL U14 ( .A0(n4), .A1(n331), .B0(n332), .Y(n333) );
  INVX1 U15 ( .A(n328), .Y(n4) );
  INVX2 U16 ( .A(n325), .Y(n386) );
  NOR2X1 U17 ( .A(n29), .B(n494), .Y(n458) );
  OAI211X1 U18 ( .A0(n5), .A1(n37), .B0(n330), .C0(n327), .Y(n335) );
  INVX1 U19 ( .A(n326), .Y(n5) );
  INVX1 U20 ( .A(n332), .Y(n330) );
  XNOR2X1 U21 ( .A(n233), .B(n442), .Y(c[1]) );
  OAI21XL U22 ( .A0(n6), .A1(n98), .B0(n325), .Y(n175) );
  INVX1 U23 ( .A(n111), .Y(n6) );
  NAND3XL U24 ( .A(n196), .B(n191), .C(n194), .Y(n205) );
  XOR3X2 U25 ( .A(n322), .B(n496), .C(n321), .Y(n339) );
  XOR3X2 U26 ( .A(n59), .B(n60), .C(n425), .Y(n427) );
  INVX1 U27 ( .A(n383), .Y(n148) );
  XOR2X1 U28 ( .A(n129), .B(n128), .Y(n383) );
  NAND2X1 U29 ( .A(n33), .B(n109), .Y(n55) );
  NAND2X1 U30 ( .A(n107), .B(n102), .Y(n449) );
  XOR2X1 U31 ( .A(n215), .B(n181), .Y(n82) );
  XNOR3X2 U32 ( .A(n252), .B(n251), .C(n250), .Y(n7) );
  XNOR3X2 U33 ( .A(n52), .B(n53), .C(n315), .Y(n8) );
  NAND2XL U34 ( .A(b[0]), .B(n500), .Y(n9) );
  INVX1 U35 ( .A(b[0]), .Y(n10) );
  INVX1 U36 ( .A(b[12]), .Y(n11) );
  INVX1 U37 ( .A(n11), .Y(n12) );
  INVX1 U38 ( .A(n11), .Y(n13) );
  INVX1 U39 ( .A(n397), .Y(n14) );
  INVX1 U40 ( .A(n224), .Y(n15) );
  NAND2BX2 U41 ( .AN(n110), .B(n111), .Y(n325) );
  BUFX3 U42 ( .A(a[12]), .Y(n111) );
  INVX1 U43 ( .A(a[10]), .Y(n16) );
  INVX1 U44 ( .A(n16), .Y(n17) );
  INVX1 U45 ( .A(n412), .Y(n18) );
  INVX1 U46 ( .A(a[8]), .Y(n19) );
  INVX1 U47 ( .A(n19), .Y(n20) );
  INVX1 U48 ( .A(n19), .Y(n21) );
  INVX1 U49 ( .A(a[7]), .Y(n22) );
  INVXL U50 ( .A(n22), .Y(n23) );
  INVX1 U51 ( .A(n493), .Y(n24) );
  INVX1 U52 ( .A(n477), .Y(n25) );
  INVX1 U53 ( .A(a[3]), .Y(n26) );
  INVXL U54 ( .A(n26), .Y(n27) );
  INVX1 U55 ( .A(n499), .Y(n28) );
  INVX1 U56 ( .A(a[1]), .Y(n29) );
  INVX1 U57 ( .A(n29), .Y(n30) );
  INVX1 U58 ( .A(n130), .Y(n31) );
  INVX1 U59 ( .A(b[8]), .Y(n32) );
  INVX1 U60 ( .A(n32), .Y(n33) );
  INVX1 U61 ( .A(n237), .Y(n34) );
  BUFX3 U62 ( .A(n110), .Y(n35) );
  INVX1 U63 ( .A(n327), .Y(n36) );
  INVX1 U64 ( .A(b[9]), .Y(n37) );
  INVX1 U65 ( .A(n37), .Y(n38) );
  INVX1 U66 ( .A(n37), .Y(n39) );
  XNOR3X4 U67 ( .A(n179), .B(n50), .C(n51), .Y(n291) );
  XOR2X2 U68 ( .A(n290), .B(n79), .Y(n297) );
  XOR2X2 U69 ( .A(n213), .B(n212), .Y(n290) );
  NAND2BX2 U70 ( .AN(n111), .B(n110), .Y(n385) );
  INVX1 U71 ( .A(b[1]), .Y(n47) );
  NAND2XL U72 ( .A(b[1]), .B(n501), .Y(n49) );
  BUFX3 U73 ( .A(a[11]), .Y(n110) );
  NOR2BX1 U74 ( .AN(n111), .B(n33), .Y(n262) );
  XOR2XL U75 ( .A(n301), .B(n8), .Y(n367) );
  XNOR3X2 U76 ( .A(n168), .B(n449), .C(n84), .Y(n50) );
  XNOR3X2 U77 ( .A(n178), .B(n177), .C(n176), .Y(n51) );
  NAND2X1 U78 ( .A(n203), .B(n202), .Y(n204) );
  XOR2X1 U79 ( .A(n82), .B(n450), .Y(c[2]) );
  NAND2XL U80 ( .A(n106), .B(n102), .Y(n440) );
  AOI22XL U81 ( .A0(n28), .A1(n457), .B0(n27), .B1(n456), .Y(n459) );
  AOI22XL U82 ( .A0(n21), .A1(n503), .B0(n18), .B1(n502), .Y(n505) );
  NAND2XL U83 ( .A(n101), .B(n108), .Y(n399) );
  AOI22XL U84 ( .A0(n17), .A1(n405), .B0(n18), .B1(n404), .Y(n406) );
  NAND2XL U85 ( .A(n96), .B(n149), .Y(n152) );
  NAND2XL U86 ( .A(n98), .B(n24), .Y(n407) );
  NAND2XL U87 ( .A(b[8]), .B(a[10]), .Y(n248) );
  NAND2XL U88 ( .A(n39), .B(n17), .Y(n266) );
  NAND2BXL U89 ( .AN(n100), .B(n111), .Y(n225) );
  NAND2XL U90 ( .A(n109), .B(n12), .Y(n324) );
  NAND2XL U91 ( .A(n101), .B(n20), .Y(n170) );
  NAND2XL U92 ( .A(n100), .B(n109), .Y(n169) );
  NAND2XL U93 ( .A(n13), .B(n105), .Y(n163) );
  NAND2XL U94 ( .A(a[3]), .B(n103), .Y(n162) );
  NAND2XL U95 ( .A(n107), .B(b[8]), .Y(n402) );
  AOI22XL U96 ( .A0(n23), .A1(n492), .B0(n21), .B1(n491), .Y(n496) );
  AOI22XL U97 ( .A0(n17), .A1(n411), .B0(n35), .B1(n410), .Y(n414) );
  INVXL U98 ( .A(n100), .Y(n237) );
  NOR2X1 U99 ( .A(n246), .B(n240), .Y(n251) );
  AOI21XL U100 ( .A0(n96), .A1(n239), .B0(n397), .Y(n240) );
  NAND2XL U101 ( .A(b[3]), .B(n21), .Y(n416) );
  INVXL U102 ( .A(n109), .Y(n412) );
  NAND2XL U103 ( .A(n17), .B(n102), .Y(n52) );
  XNOR2X1 U104 ( .A(n303), .B(n302), .Y(n53) );
  NAND2XL U105 ( .A(a[12]), .B(n13), .Y(n371) );
  NAND2XL U106 ( .A(n23), .B(n13), .Y(n286) );
  NAND2XL U107 ( .A(n96), .B(n304), .Y(n314) );
  NAND2XL U108 ( .A(a[7]), .B(n31), .Y(n247) );
  NAND2XL U109 ( .A(n108), .B(n36), .Y(n451) );
  NAND2XL U110 ( .A(n38), .B(n109), .Y(n249) );
  NAND2XL U111 ( .A(n27), .B(b[4]), .Y(n489) );
  NAND2XL U112 ( .A(b[4]), .B(n30), .Y(n470) );
  INVXL U113 ( .A(n101), .Y(n397) );
  NAND2XL U114 ( .A(n107), .B(n13), .Y(n222) );
  NAND2XL U115 ( .A(n100), .B(n108), .Y(n418) );
  NAND2XL U116 ( .A(n108), .B(n33), .Y(n438) );
  NAND2XL U117 ( .A(n107), .B(n38), .Y(n441) );
  NAND2XL U118 ( .A(n97), .B(n18), .Y(n422) );
  NAND2XL U119 ( .A(n98), .B(n21), .Y(n421) );
  NAND2XL U120 ( .A(a[7]), .B(n102), .Y(n465) );
  NAND2XL U121 ( .A(n109), .B(n103), .Y(n302) );
  NAND2XL U122 ( .A(n21), .B(n31), .Y(n280) );
  NAND2XL U123 ( .A(n108), .B(n12), .Y(n235) );
  NAND2XL U124 ( .A(a[7]), .B(b[8]), .Y(n448) );
  NAND2XL U125 ( .A(n100), .B(n104), .Y(n472) );
  NAND2XL U126 ( .A(n101), .B(a[10]), .Y(n223) );
  NAND2XL U127 ( .A(n20), .B(n102), .Y(n236) );
  NAND2XL U128 ( .A(n108), .B(n103), .Y(n464) );
  NAND2XL U129 ( .A(n104), .B(n31), .Y(n372) );
  NAND2XL U130 ( .A(n20), .B(n12), .Y(n303) );
  INVXL U131 ( .A(n107), .Y(n395) );
  NAND2XL U132 ( .A(n96), .B(n261), .Y(n264) );
  XNOR3X2 U133 ( .A(n54), .B(n55), .C(n228), .Y(n230) );
  NAND2XL U134 ( .A(n38), .B(n21), .Y(n54) );
  NAND2XL U135 ( .A(n101), .B(a[7]), .Y(n439) );
  NAND2XL U136 ( .A(n100), .B(a[7]), .Y(n400) );
  NAND2XL U137 ( .A(n100), .B(n17), .Y(n187) );
  NAND2XL U138 ( .A(a[5]), .B(b[3]), .Y(n498) );
  NAND2XL U139 ( .A(n101), .B(n27), .Y(n362) );
  NAND2XL U140 ( .A(n107), .B(n99), .Y(n361) );
  NAND2BXL U141 ( .AN(n100), .B(n110), .Y(n239) );
  NAND2XL U142 ( .A(a[3]), .B(n97), .Y(n481) );
  NAND2XL U143 ( .A(n105), .B(n98), .Y(n480) );
  XOR3X2 U144 ( .A(n57), .B(n415), .C(n373), .Y(n374) );
  NAND2XL U145 ( .A(a[1]), .B(n36), .Y(n57) );
  XOR3X2 U146 ( .A(n58), .B(n316), .C(n367), .Y(n317) );
  NAND2XL U147 ( .A(n34), .B(n30), .Y(n58) );
  XNOR3X2 U148 ( .A(n417), .B(n384), .C(n383), .Y(n59) );
  XNOR2X1 U149 ( .A(n419), .B(n418), .Y(n60) );
  NAND2XL U150 ( .A(a[0]), .B(n13), .Y(n426) );
  XOR3X2 U151 ( .A(n61), .B(n497), .C(n376), .Y(n337) );
  NAND2XL U152 ( .A(n104), .B(n33), .Y(n61) );
  XOR3X2 U153 ( .A(n62), .B(n360), .C(n359), .Y(n364) );
  NAND2XL U154 ( .A(n21), .B(b[2]), .Y(n62) );
  XOR3X2 U155 ( .A(n63), .B(n409), .C(n95), .Y(n375) );
  NAND2XL U156 ( .A(a[3]), .B(n33), .Y(n63) );
  NAND2XL U157 ( .A(n13), .B(a[1]), .Y(n141) );
  NAND2XL U158 ( .A(n103), .B(n105), .Y(n142) );
  NAND2XL U159 ( .A(n102), .B(a[3]), .Y(n143) );
  NAND2XL U160 ( .A(n100), .B(n20), .Y(n87) );
  NAND2XL U161 ( .A(n109), .B(n99), .Y(n92) );
  NAND2XL U162 ( .A(n21), .B(n99), .Y(n85) );
  NAND2XL U163 ( .A(n109), .B(n98), .Y(n86) );
  NAND2XL U164 ( .A(n33), .B(n30), .Y(n353) );
  NAND2BXL U165 ( .AN(b[2]), .B(n110), .Y(n149) );
  NAND2BXL U166 ( .AN(b[8]), .B(n35), .Y(n304) );
  NAND2BXL U167 ( .AN(n101), .B(n35), .Y(n261) );
  BUFX8 U168 ( .A(n385), .Y(n96) );
  OAI2BB1X1 U169 ( .A0N(n110), .A1N(n327), .B0(n96), .Y(n127) );
  AOI22XL U170 ( .A0(n27), .A1(n461), .B0(n106), .B1(n460), .Y(n463) );
  NAND2XL U171 ( .A(n106), .B(n13), .Y(n453) );
  NAND2XL U172 ( .A(n107), .B(n103), .Y(n454) );
  AND2X1 U173 ( .A(n106), .B(n103), .Y(n84) );
  AND2X1 U174 ( .A(n17), .B(n98), .Y(n155) );
  AND2X1 U175 ( .A(n17), .B(n97), .Y(n140) );
  AND2X1 U176 ( .A(n109), .B(n102), .Y(n278) );
  AND2X1 U177 ( .A(n34), .B(n105), .Y(n322) );
  AND2X1 U178 ( .A(n104), .B(n98), .Y(n220) );
  INVXL U179 ( .A(n103), .Y(n130) );
  NAND2XL U180 ( .A(n14), .B(n105), .Y(n350) );
  NAND2XL U181 ( .A(n107), .B(n34), .Y(n369) );
  NAND2XL U182 ( .A(n34), .B(n27), .Y(n349) );
  NAND2XL U183 ( .A(b[4]), .B(a[5]), .Y(n506) );
  NAND2XL U184 ( .A(n25), .B(n34), .Y(n357) );
  NAND2XL U185 ( .A(n14), .B(n30), .Y(n319) );
  NAND2XL U186 ( .A(n27), .B(b[2]), .Y(n469) );
  NAND2XL U187 ( .A(n33), .B(n105), .Y(n358) );
  NAND2XL U188 ( .A(n15), .B(n27), .Y(n320) );
  NAND2XL U189 ( .A(n25), .B(n14), .Y(n368) );
  NAND2XL U190 ( .A(n28), .B(n36), .Y(n431) );
  NAND2XL U191 ( .A(n30), .B(n31), .Y(n430) );
  NAND2XL U192 ( .A(n25), .B(n33), .Y(n429) );
  NAND2XL U193 ( .A(n27), .B(n39), .Y(n428) );
  NAND2XL U194 ( .A(b[1]), .B(n501), .Y(n65) );
  OAI2BB1X1 U195 ( .A0N(b[2]), .A1N(n137), .B0(n136), .Y(n139) );
  NAND2XL U196 ( .A(n96), .B(n134), .Y(n137) );
  NAND2BXL U197 ( .AN(b[1]), .B(n35), .Y(n134) );
  NAND2XL U198 ( .A(b[2]), .B(n17), .Y(n420) );
  AOI2BB2XL U199 ( .B0(b[0]), .B1(n386), .A0N(n96), .A1N(n500), .Y(n387) );
  NAND2XL U200 ( .A(b[0]), .B(n500), .Y(n66) );
  XNOR2X1 U201 ( .A(n148), .B(n180), .Y(n366) );
  XNOR2X1 U202 ( .A(n79), .B(n7), .Y(n321) );
  XOR2X1 U203 ( .A(n148), .B(n384), .Y(n67) );
  XOR3X2 U204 ( .A(n367), .B(n366), .C(n365), .Y(c[10]) );
  NAND3X1 U205 ( .A(n64), .B(n330), .C(n328), .Y(n334) );
  XOR2X1 U206 ( .A(n447), .B(n448), .Y(n179) );
  XNOR3X2 U207 ( .A(n67), .B(n181), .C(n214), .Y(n233) );
  NOR2X1 U208 ( .A(n64), .B(n327), .Y(n331) );
  XOR3X2 U209 ( .A(n215), .B(n290), .C(n214), .Y(n216) );
  XNOR3X2 U210 ( .A(n382), .B(n381), .C(n380), .Y(c[11]) );
  XNOR3X2 U211 ( .A(n370), .B(n369), .C(n368), .Y(n382) );
  XOR2X1 U212 ( .A(n375), .B(n374), .Y(n381) );
  XNOR3X2 U213 ( .A(n378), .B(n377), .C(n376), .Y(n380) );
  XNOR3X2 U214 ( .A(n321), .B(n82), .C(n260), .Y(c[5]) );
  XNOR3X2 U215 ( .A(n468), .B(n259), .C(n254), .Y(n260) );
  XOR2X1 U216 ( .A(n253), .B(n469), .Y(n254) );
  XNOR2X1 U217 ( .A(n471), .B(n470), .Y(n259) );
  XNOR3X2 U218 ( .A(n343), .B(n339), .C(n338), .Y(c[8]) );
  XOR2X1 U219 ( .A(n320), .B(n319), .Y(n343) );
  XNOR2X1 U220 ( .A(n337), .B(n336), .Y(n338) );
  INVX1 U221 ( .A(n371), .Y(n384) );
  NOR2X1 U222 ( .A(n395), .B(n397), .Y(n417) );
  XOR3X2 U223 ( .A(n68), .B(n77), .C(n78), .Y(n365) );
  XNOR3X2 U224 ( .A(n408), .B(n407), .C(n406), .Y(n68) );
  XOR2X1 U225 ( .A(n358), .B(n357), .Y(n77) );
  XNOR2X1 U226 ( .A(n364), .B(n363), .Y(n78) );
  XOR2X1 U227 ( .A(n236), .B(n235), .Y(n252) );
  XOR3X2 U228 ( .A(n249), .B(n248), .C(n247), .Y(n250) );
  NAND2XL U229 ( .A(n202), .B(n195), .Y(n210) );
  INVX1 U230 ( .A(n373), .Y(n180) );
  XOR3X2 U231 ( .A(n80), .B(n81), .C(n230), .Y(n79) );
  XNOR2X1 U232 ( .A(n223), .B(n222), .Y(n80) );
  XOR2X1 U233 ( .A(n464), .B(n465), .Y(n81) );
  XOR2X1 U234 ( .A(n394), .B(n8), .Y(n376) );
  XNOR3X2 U235 ( .A(n83), .B(n296), .C(n292), .Y(c[6]) );
  XNOR3X2 U236 ( .A(n384), .B(n291), .C(n290), .Y(n292) );
  XOR2X1 U237 ( .A(n435), .B(n434), .Y(c[12]) );
  XOR2X1 U238 ( .A(n433), .B(n432), .Y(n434) );
  INVX1 U239 ( .A(n196), .Y(n202) );
  INVX1 U240 ( .A(n385), .Y(n192) );
  XNOR2X1 U241 ( .A(n301), .B(n7), .Y(n83) );
  XOR2X1 U242 ( .A(n318), .B(n317), .Y(c[7]) );
  XOR2X1 U243 ( .A(n217), .B(n216), .Y(c[3]) );
  XNOR3X2 U244 ( .A(n83), .B(n356), .C(n355), .Y(c[9]) );
  NOR2XL U245 ( .A(n494), .B(n395), .Y(n487) );
  OAI21XL U246 ( .A0(n18), .A1(n47), .B0(n49), .Y(n503) );
  OAI21XL U247 ( .A0(n21), .A1(n501), .B0(n66), .Y(n502) );
  OAI21XL U248 ( .A0(n27), .A1(n47), .B0(n49), .Y(n457) );
  OAI21XL U249 ( .A0(n105), .A1(n501), .B0(n66), .Y(n456) );
  OAI21XL U250 ( .A0(n17), .A1(n47), .B0(n49), .Y(n404) );
  OAI21XL U251 ( .A0(n18), .A1(n501), .B0(n9), .Y(n405) );
  OAI21XL U252 ( .A0(a[5]), .A1(n47), .B0(n49), .Y(n467) );
  OAI21XL U253 ( .A0(n106), .A1(n501), .B0(n9), .Y(n466) );
  OAI21XL U254 ( .A0(n108), .A1(n500), .B0(n65), .Y(n476) );
  OAI21XL U255 ( .A0(n106), .A1(n47), .B0(n49), .Y(n461) );
  OAI21XL U256 ( .A0(n107), .A1(n501), .B0(n9), .Y(n475) );
  OAI21XL U257 ( .A0(n30), .A1(n10), .B0(n66), .Y(n443) );
  OAI21XL U258 ( .A0(n27), .A1(n501), .B0(n9), .Y(n460) );
  OAI21XL U259 ( .A0(n24), .A1(n10), .B0(n66), .Y(n485) );
  XNOR3X2 U260 ( .A(n440), .B(n165), .C(n164), .Y(n166) );
  XNOR3X2 U261 ( .A(n155), .B(n154), .C(n153), .Y(n167) );
  INVX1 U262 ( .A(b[2]), .Y(n494) );
  NAND2X1 U263 ( .A(n39), .B(n326), .Y(n328) );
  XNOR3X2 U264 ( .A(n451), .B(n452), .C(n211), .Y(n212) );
  NAND3X1 U265 ( .A(n210), .B(n205), .C(n204), .Y(n213) );
  NAND2X1 U266 ( .A(n23), .B(n39), .Y(n452) );
  XOR3X2 U267 ( .A(n189), .B(n188), .C(n187), .Y(n196) );
  NAND2X1 U268 ( .A(b[8]), .B(n20), .Y(n188) );
  NAND2X1 U269 ( .A(n101), .B(n109), .Y(n189) );
  XOR2X1 U270 ( .A(n289), .B(n288), .Y(n301) );
  XOR2X1 U271 ( .A(n286), .B(n280), .Y(n288) );
  XNOR3X2 U272 ( .A(n278), .B(n266), .C(n265), .Y(n289) );
  OAI2BB1X1 U273 ( .A0N(n13), .A1N(n133), .B0(n132), .Y(n373) );
  OAI21XL U274 ( .A0(n131), .A1(n386), .B0(n31), .Y(n132) );
  OAI2BB1X1 U275 ( .A0N(n35), .A1N(n130), .B0(n96), .Y(n133) );
  NOR2BX1 U276 ( .AN(a[12]), .B(n13), .Y(n131) );
  NOR2BX1 U277 ( .AN(n111), .B(n103), .Y(n122) );
  NOR2BX1 U278 ( .AN(n110), .B(n97), .Y(n173) );
  XNOR2X1 U279 ( .A(n324), .B(n323), .Y(n332) );
  NAND2X1 U280 ( .A(a[10]), .B(n103), .Y(n323) );
  XOR2X1 U281 ( .A(n147), .B(n146), .Y(n214) );
  XNOR3X2 U282 ( .A(n399), .B(n145), .C(n144), .Y(n146) );
  XNOR3X2 U283 ( .A(n140), .B(n139), .C(n138), .Y(n147) );
  XNOR3X2 U284 ( .A(n383), .B(n348), .C(n347), .Y(n356) );
  XOR2X1 U285 ( .A(n346), .B(n506), .Y(n347) );
  XNOR2X1 U286 ( .A(n507), .B(n504), .Y(n348) );
  NAND2X1 U287 ( .A(n25), .B(n15), .Y(n346) );
  NAND2X1 U288 ( .A(b[4]), .B(n23), .Y(n415) );
  XOR2X1 U289 ( .A(n300), .B(n299), .Y(n316) );
  NAND2X1 U290 ( .A(n104), .B(n14), .Y(n299) );
  XNOR3X2 U291 ( .A(n234), .B(n297), .C(n233), .Y(c[4]) );
  XOR2X1 U292 ( .A(n463), .B(n221), .Y(n234) );
  XOR3X2 U293 ( .A(n220), .B(n219), .C(n462), .Y(n221) );
  XOR2X1 U294 ( .A(n170), .B(n169), .Y(n177) );
  XOR2X1 U295 ( .A(n163), .B(n162), .Y(n165) );
  XOR2X1 U296 ( .A(n401), .B(n402), .Y(n145) );
  NAND2X1 U297 ( .A(n106), .B(n38), .Y(n401) );
  XOR3X2 U298 ( .A(n426), .B(n427), .C(n394), .Y(n435) );
  XOR2X1 U299 ( .A(n424), .B(n423), .Y(n425) );
  XNOR3X2 U300 ( .A(n488), .B(n298), .C(n297), .Y(n318) );
  XOR3X2 U301 ( .A(n489), .B(n490), .C(n487), .Y(n298) );
  AOI22X1 U302 ( .A0(n24), .A1(n486), .B0(n23), .B1(n485), .Y(n488) );
  NAND2X1 U303 ( .A(n106), .B(b[3]), .Y(n490) );
  XNOR3X2 U304 ( .A(n67), .B(n455), .C(n182), .Y(n217) );
  NOR2X1 U305 ( .A(n396), .B(n398), .Y(n455) );
  XNOR2X1 U306 ( .A(n458), .B(n459), .Y(n182) );
  INVX1 U307 ( .A(n97), .Y(n398) );
  XOR2X1 U308 ( .A(n422), .B(n421), .Y(n423) );
  XOR2X1 U309 ( .A(n481), .B(n480), .Y(n482) );
  NAND2X1 U310 ( .A(n106), .B(b[4]), .Y(n497) );
  OAI2BB1X1 U311 ( .A0N(n110), .A1N(n224), .B0(n96), .Y(n227) );
  NAND2X1 U312 ( .A(n108), .B(n38), .Y(n447) );
  OAI2BB1X1 U313 ( .A0N(n97), .A1N(n175), .B0(n174), .Y(n176) );
  OAI21XL U314 ( .A0(n173), .A1(n192), .B0(n98), .Y(n174) );
  NAND2BX1 U315 ( .AN(n66), .B(a[12]), .Y(n388) );
  XNOR3X2 U316 ( .A(n85), .B(n86), .C(n400), .Y(n138) );
  XOR3X2 U317 ( .A(n143), .B(n142), .C(n141), .Y(n144) );
  XOR2X1 U318 ( .A(n446), .B(n445), .Y(n450) );
  NOR2X1 U319 ( .A(n396), .B(n494), .Y(n445) );
  AOI22X1 U320 ( .A0(n30), .A1(n444), .B0(n28), .B1(n443), .Y(n446) );
  OAI21XL U321 ( .A0(n28), .A1(n47), .B0(n49), .Y(n444) );
  XNOR3X2 U322 ( .A(n354), .B(n353), .C(n352), .Y(n355) );
  XOR3X2 U323 ( .A(n351), .B(n350), .C(n349), .Y(n352) );
  XOR2X1 U324 ( .A(n394), .B(n505), .Y(n354) );
  AOI21X1 U325 ( .A0(n100), .A1(n227), .B0(n226), .Y(n228) );
  OAI2BB1X1 U326 ( .A0N(n33), .A1N(n264), .B0(n263), .Y(n265) );
  OAI21XL U327 ( .A0(n262), .A1(n386), .B0(n101), .Y(n263) );
  XNOR3X2 U328 ( .A(n403), .B(n366), .C(n214), .Y(c[0]) );
  NOR2X1 U329 ( .A(n396), .B(n10), .Y(n403) );
  XOR2X1 U330 ( .A(n479), .B(n478), .Y(n483) );
  NOR2X1 U331 ( .A(n494), .B(n477), .Y(n478) );
  AOI22X1 U332 ( .A0(n107), .A1(n476), .B0(n108), .B1(n475), .Y(n479) );
  INVX1 U333 ( .A(n106), .Y(n477) );
  NAND2X1 U334 ( .A(n99), .B(n23), .Y(n419) );
  XOR2X1 U335 ( .A(n484), .B(n474), .Y(n296) );
  XOR2X1 U336 ( .A(n473), .B(n472), .Y(n474) );
  XOR2X1 U337 ( .A(n483), .B(n482), .Y(n484) );
  NAND2X1 U338 ( .A(n99), .B(a[1]), .Y(n473) );
  INVX1 U339 ( .A(n191), .Y(n195) );
  OAI21XL U340 ( .A0(n190), .A1(n386), .B0(n98), .Y(n191) );
  NOR2BX1 U341 ( .AN(a[12]), .B(n99), .Y(n190) );
  INVX1 U342 ( .A(n194), .Y(n203) );
  OAI21XL U343 ( .A0(n193), .A1(n192), .B0(n99), .Y(n194) );
  NOR2BX1 U344 ( .AN(n110), .B(n98), .Y(n193) );
  OAI21XL U345 ( .A0(n21), .A1(n47), .B0(n49), .Y(n492) );
  OAI21XL U346 ( .A0(n23), .A1(n501), .B0(n66), .Y(n491) );
  INVX1 U347 ( .A(n414), .Y(n377) );
  OAI21XL U348 ( .A0(n35), .A1(n47), .B0(n49), .Y(n411) );
  OAI21XL U349 ( .A0(n17), .A1(n501), .B0(n9), .Y(n410) );
  NAND2BXL U350 ( .AN(n101), .B(n111), .Y(n238) );
  OAI2BB1X1 U351 ( .A0N(n39), .A1N(n314), .B0(n306), .Y(n315) );
  OAI21XL U352 ( .A0(n305), .A1(n386), .B0(n33), .Y(n306) );
  NOR2BX1 U353 ( .AN(n111), .B(n39), .Y(n305) );
  OAI2BB1X1 U354 ( .A0N(n97), .A1N(n152), .B0(n151), .Y(n154) );
  OAI21XL U355 ( .A0(n150), .A1(n386), .B0(b[2]), .Y(n151) );
  NOR2BX1 U356 ( .AN(n111), .B(n97), .Y(n150) );
  AND2X2 U357 ( .A(n12), .B(a[3]), .Y(n168) );
  XNOR3X2 U358 ( .A(n87), .B(n92), .C(n439), .Y(n153) );
  AND2X2 U359 ( .A(a[10]), .B(n99), .Y(n178) );
  XNOR2X1 U360 ( .A(n441), .B(n438), .Y(n164) );
  XNOR2X1 U361 ( .A(n453), .B(n454), .Y(n211) );
  INVX1 U362 ( .A(n102), .Y(n327) );
  INVX1 U363 ( .A(n99), .Y(n224) );
  OAI21XL U364 ( .A0(n23), .A1(n47), .B0(n49), .Y(n486) );
  NOR2X1 U365 ( .A(n494), .B(n499), .Y(n462) );
  INVX1 U366 ( .A(n105), .Y(n499) );
  NAND2X1 U367 ( .A(n105), .B(n39), .Y(n409) );
  XOR2X1 U368 ( .A(n372), .B(n371), .Y(n95) );
  NAND2X1 U369 ( .A(n104), .B(n36), .Y(n359) );
  NAND2X1 U370 ( .A(n39), .B(a[1]), .Y(n360) );
  XOR2X1 U371 ( .A(n362), .B(n361), .Y(n363) );
  XOR2X1 U372 ( .A(n431), .B(n430), .Y(n432) );
  XOR2X1 U373 ( .A(n498), .B(n495), .Y(n336) );
  NOR2X1 U374 ( .A(n494), .B(n493), .Y(n495) );
  INVX1 U375 ( .A(n108), .Y(n493) );
  AND2X2 U376 ( .A(n97), .B(a[1]), .Y(n219) );
  NAND2X1 U377 ( .A(n15), .B(n28), .Y(n300) );
  NAND2X1 U378 ( .A(n104), .B(n15), .Y(n253) );
  NAND2X1 U379 ( .A(b[3]), .B(n24), .Y(n507) );
  NAND2X1 U380 ( .A(n105), .B(b[3]), .Y(n471) );
  AND2X2 U381 ( .A(n23), .B(b[2]), .Y(n504) );
  NAND2X1 U382 ( .A(n97), .B(n23), .Y(n408) );
  NAND2X1 U383 ( .A(n104), .B(n39), .Y(n351) );
  NAND2X1 U384 ( .A(n24), .B(n99), .Y(n370) );
  INVX1 U385 ( .A(n104), .Y(n396) );
  XOR2X1 U386 ( .A(n429), .B(n428), .Y(n433) );
  AOI22X1 U387 ( .A0(a[0]), .A1(n437), .B0(n30), .B1(n436), .Y(n442) );
  OAI21XL U388 ( .A0(n30), .A1(n47), .B0(n49), .Y(n437) );
  OAI21XL U389 ( .A0(n104), .A1(n10), .B0(n9), .Y(n436) );
  XOR2X1 U390 ( .A(n416), .B(n413), .Y(n378) );
  NOR2X1 U391 ( .A(n412), .B(n494), .Y(n413) );
  INVX1 U392 ( .A(b[0]), .Y(n501) );
  INVX1 U393 ( .A(b[1]), .Y(n500) );
  BUFX3 U394 ( .A(a[4]), .Y(n106) );
  BUFX3 U395 ( .A(a[6]), .Y(n108) );
  BUFX3 U396 ( .A(a[2]), .Y(n105) );
  BUFX3 U397 ( .A(a[5]), .Y(n107) );
  BUFX3 U398 ( .A(b[11]), .Y(n103) );
  BUFX3 U399 ( .A(a[9]), .Y(n109) );
  BUFX3 U400 ( .A(b[10]), .Y(n102) );
  BUFX3 U401 ( .A(b[4]), .Y(n98) );
  BUFX3 U402 ( .A(b[7]), .Y(n101) );
  BUFX3 U403 ( .A(b[3]), .Y(n97) );
  BUFX3 U404 ( .A(b[5]), .Y(n99) );
  BUFX3 U405 ( .A(b[6]), .Y(n100) );
  BUFX3 U406 ( .A(a[0]), .Y(n104) );
  XOR2X1 U407 ( .A(n389), .B(n420), .Y(n424) );
  OAI21XL U408 ( .A0(n135), .A1(n386), .B0(b[1]), .Y(n136) );
  NOR2BX1 U409 ( .AN(a[12]), .B(b[2]), .Y(n135) );
  AOI21XL U410 ( .A0(n325), .A1(n238), .B0(n237), .Y(n246) );
  AOI21XL U411 ( .A0(n325), .A1(n225), .B0(n224), .Y(n226) );
endmodule


module multiplier_12 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n36, n37, n38, n39, n43, n47, n49, n50, n51, n52,
         n53, n54, n55, n57, n58, n59, n61, n63, n64, n77, n81, n83, n84, n85,
         n86, n87, n92, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n122, n127, n128, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n202, n203, n204, n205, n210,
         n211, n212, n213, n214, n215, n216, n217, n219, n220, n221, n239,
         n240, n246, n247, n248, n249, n250, n251, n252, n253, n254, n259,
         n260, n261, n262, n263, n264, n265, n266, n286, n288, n289, n290,
         n291, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n311, n314, n315, n316, n317, n318, n319, n320, n321, n323,
         n324, n325, n326, n327, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538;

  BUFX4 U1 ( .A(b[5]), .Y(n96) );
  XOR2X2 U2 ( .A(n249), .B(n248), .Y(n296) );
  OAI21X1 U3 ( .A0(n374), .A1(n373), .B0(n372), .Y(n448) );
  AND2X2 U4 ( .A(n169), .B(n92), .Y(n371) );
  AOI211X1 U5 ( .A0(n96), .A1(n37), .B0(n34), .C0(n170), .Y(n1) );
  INVX1 U6 ( .A(n1), .Y(n173) );
  NOR2X1 U7 ( .A(n31), .B(n34), .Y(n300) );
  OAI21XL U8 ( .A0(n98), .A1(n365), .B0(n367), .Y(n220) );
  NAND2XL U9 ( .A(n25), .B(n92), .Y(n537) );
  OAI221XL U10 ( .A0(n34), .A1(n7), .B0(n365), .B1(n59), .C0(n368), .Y(n369)
         );
  NOR2XL U11 ( .A(n385), .B(n388), .Y(n470) );
  NAND2X1 U12 ( .A(n30), .B(n14), .Y(n239) );
  NAND2XL U13 ( .A(n24), .B(n92), .Y(n405) );
  NOR2X1 U14 ( .A(n5), .B(n34), .Y(n217) );
  NOR2X1 U15 ( .A(n31), .B(n365), .Y(n315) );
  NOR2XL U16 ( .A(n519), .B(n16), .Y(n411) );
  INVX1 U17 ( .A(n92), .Y(n388) );
  XOR3X2 U18 ( .A(n350), .B(n334), .C(n349), .Y(c[10]) );
  XNOR3X2 U19 ( .A(n376), .B(n465), .C(n181), .Y(c[2]) );
  OAI2BB1XL U20 ( .A0N(n36), .A1N(n314), .B0(n311), .Y(n317) );
  AOI21XL U21 ( .A0(n311), .A1(n253), .B0(n252), .Y(n260) );
  AOI21XL U22 ( .A0(n311), .A1(n189), .B0(n188), .Y(n190) );
  XNOR3X2 U23 ( .A(n210), .B(n205), .C(n204), .Y(n382) );
  AOI21X1 U24 ( .A0(n97), .A1(n191), .B0(n190), .Y(n210) );
  NAND2BX1 U25 ( .AN(a[11]), .B(a[12]), .Y(n311) );
  INVX1 U26 ( .A(n492), .Y(n381) );
  XOR2X2 U27 ( .A(n165), .B(n164), .Y(n376) );
  NAND2XL U28 ( .A(n4), .B(n20), .Y(n168) );
  NAND2X1 U29 ( .A(n18), .B(b[11]), .Y(n297) );
  XOR2X2 U30 ( .A(n47), .B(n178), .Y(n43) );
  MXI2X1 U31 ( .A(n34), .B(n371), .S0(n95), .Y(n374) );
  BUFX3 U32 ( .A(n367), .Y(n86) );
  NAND2BX1 U33 ( .AN(a[12]), .B(a[11]), .Y(n367) );
  NAND2BX1 U34 ( .AN(a[12]), .B(a[11]), .Y(n169) );
  XOR2X1 U35 ( .A(n464), .B(n463), .Y(n492) );
  AOI21X2 U36 ( .A0(n33), .A1(n110), .B0(n109), .Y(n111) );
  XOR2X1 U37 ( .A(n538), .B(n2), .Y(n352) );
  INVX1 U38 ( .A(n34), .Y(n36) );
  INVX1 U39 ( .A(n99), .Y(n314) );
  INVX1 U40 ( .A(a[11]), .Y(n365) );
  INVX1 U41 ( .A(a[12]), .Y(n34) );
  XNOR3X2 U42 ( .A(n55), .B(n57), .C(n303), .Y(n2) );
  INVX1 U43 ( .A(b[8]), .Y(n3) );
  INVX1 U44 ( .A(n3), .Y(n4) );
  INVX1 U45 ( .A(n3), .Y(n5) );
  INVX1 U46 ( .A(n387), .Y(n6) );
  NAND2XL U47 ( .A(b[0]), .B(n531), .Y(n7) );
  NAND2X1 U48 ( .A(b[0]), .B(n531), .Y(n58) );
  BUFX3 U49 ( .A(n59), .Y(n8) );
  NAND2X1 U50 ( .A(b[1]), .B(n532), .Y(n59) );
  INVX1 U51 ( .A(b[0]), .Y(n9) );
  INVX1 U52 ( .A(n188), .Y(n10) );
  BUFX3 U53 ( .A(n92), .Y(n11) );
  BUFX3 U54 ( .A(b[3]), .Y(n92) );
  INVX1 U55 ( .A(n386), .Y(n12) );
  INVX1 U56 ( .A(a[10]), .Y(n13) );
  INVX1 U57 ( .A(n13), .Y(n14) );
  INVX1 U58 ( .A(n13), .Y(n15) );
  INVX1 U59 ( .A(a[9]), .Y(n16) );
  INVX1 U60 ( .A(n16), .Y(n17) );
  INVX1 U61 ( .A(n16), .Y(n18) );
  INVX1 U62 ( .A(a[8]), .Y(n19) );
  INVX1 U63 ( .A(n19), .Y(n20) );
  INVX1 U64 ( .A(n19), .Y(n21) );
  INVX1 U65 ( .A(a[7]), .Y(n22) );
  INVX1 U66 ( .A(n22), .Y(n23) );
  INVXL U67 ( .A(n22), .Y(n24) );
  INVX1 U68 ( .A(n518), .Y(n25) );
  INVX1 U69 ( .A(n498), .Y(n26) );
  INVX1 U70 ( .A(n462), .Y(n27) );
  NAND2X1 U71 ( .A(n104), .B(b[11]), .Y(n152) );
  INVX1 U72 ( .A(n530), .Y(n28) );
  INVX1 U73 ( .A(b[9]), .Y(n29) );
  INVX1 U74 ( .A(n29), .Y(n30) );
  INVX1 U75 ( .A(n29), .Y(n31) );
  INVX1 U76 ( .A(n252), .Y(n32) );
  BUFX3 U77 ( .A(b[6]), .Y(n97) );
  BUFX3 U78 ( .A(b[4]), .Y(n95) );
  AOI21X1 U79 ( .A0(n311), .A1(n108), .B0(n314), .Y(n109) );
  INVX1 U80 ( .A(n311), .Y(n373) );
  AOI22X1 U81 ( .A0(n12), .A1(n127), .B0(n33), .B1(n122), .Y(n377) );
  NOR2X2 U82 ( .A(n260), .B(n259), .Y(n265) );
  AOI21XL U83 ( .A0(n86), .A1(n254), .B0(n387), .Y(n259) );
  XOR2X2 U84 ( .A(n143), .B(n142), .Y(n179) );
  OAI21XL U85 ( .A0(n15), .A1(n366), .B0(n59), .Y(n400) );
  OAI21XL U86 ( .A0(n107), .A1(n366), .B0(n59), .Y(n497) );
  XNOR3X4 U87 ( .A(n377), .B(n53), .C(n376), .Y(n378) );
  BUFX3 U88 ( .A(b[11]), .Y(n33) );
  NAND2XL U89 ( .A(n107), .B(n33), .Y(n480) );
  NAND2XL U90 ( .A(n99), .B(n104), .Y(n132) );
  BUFX3 U91 ( .A(b[10]), .Y(n99) );
  NOR2BXL U92 ( .AN(a[12]), .B(n92), .Y(n146) );
  INVX1 U93 ( .A(n365), .Y(n37) );
  OAI2BB1X4 U94 ( .A0N(a[11]), .A1N(n314), .B0(n86), .Y(n110) );
  INVX2 U95 ( .A(n144), .Y(n330) );
  INVXL U96 ( .A(n288), .Y(n215) );
  NAND2X1 U97 ( .A(n98), .B(n17), .Y(n167) );
  INVX1 U98 ( .A(n96), .Y(n188) );
  XOR2X1 U99 ( .A(n491), .B(n490), .Y(c[5]) );
  XNOR3X2 U100 ( .A(n363), .B(n362), .C(n361), .Y(c[11]) );
  NAND2XL U101 ( .A(n106), .B(n33), .Y(n469) );
  NAND2XL U102 ( .A(n104), .B(n92), .Y(n502) );
  NAND2XL U103 ( .A(n105), .B(n11), .Y(n511) );
  INVXL U104 ( .A(n364), .Y(n180) );
  XOR3X2 U105 ( .A(n39), .B(n265), .C(n264), .Y(n38) );
  XNOR2X1 U106 ( .A(n251), .B(n250), .Y(n39) );
  XOR3X2 U107 ( .A(n466), .B(n467), .C(n166), .Y(n47) );
  NOR2XL U108 ( .A(n383), .B(n387), .Y(n415) );
  XOR2XL U109 ( .A(n296), .B(n2), .Y(n334) );
  NOR2XL U110 ( .A(n384), .B(n387), .Y(n512) );
  XNOR2X1 U111 ( .A(n492), .B(n377), .Y(n181) );
  XOR3X2 U112 ( .A(n49), .B(n402), .C(n50), .Y(n349) );
  XOR3X2 U113 ( .A(n403), .B(n336), .C(n335), .Y(n49) );
  XNOR3X2 U114 ( .A(n348), .B(n347), .C(n346), .Y(n50) );
  XNOR2X1 U115 ( .A(n330), .B(n64), .Y(n364) );
  XOR2X1 U116 ( .A(n63), .B(n443), .Y(c[1]) );
  NAND2XL U117 ( .A(n98), .B(n107), .Y(n395) );
  NAND2XL U118 ( .A(n6), .B(n104), .Y(n336) );
  NAND2XL U119 ( .A(n24), .B(n31), .Y(n467) );
  NAND2XL U120 ( .A(n98), .B(n21), .Y(n450) );
  AOI22XL U121 ( .A0(n21), .A1(n534), .B0(n18), .B1(n533), .Y(n535) );
  OAI21XL U122 ( .A0(n174), .A1(n188), .B0(n173), .Y(n175) );
  NAND2XL U123 ( .A(n105), .B(n30), .Y(n397) );
  NAND2XL U124 ( .A(n106), .B(n4), .Y(n398) );
  NAND2XL U125 ( .A(n100), .B(n103), .Y(n153) );
  NAND2BXL U126 ( .AN(n97), .B(n36), .Y(n189) );
  INVXL U127 ( .A(n98), .Y(n387) );
  NAND2XL U128 ( .A(n24), .B(n12), .Y(n247) );
  NAND2XL U129 ( .A(n21), .B(n99), .Y(n261) );
  OAI21XL U130 ( .A0(n315), .A1(n370), .B0(n99), .Y(n316) );
  XNOR3X2 U131 ( .A(n51), .B(n408), .C(n318), .Y(n538) );
  NAND2XL U132 ( .A(n18), .B(n100), .Y(n51) );
  INVX1 U133 ( .A(n169), .Y(n370) );
  OAI2BB1X1 U134 ( .A0N(n92), .A1N(n148), .B0(n147), .Y(n150) );
  NAND2XL U135 ( .A(n86), .B(n145), .Y(n148) );
  NAND2BXL U136 ( .AN(n87), .B(a[11]), .Y(n145) );
  NAND2XL U137 ( .A(n95), .B(n106), .Y(n536) );
  XNOR3X2 U138 ( .A(n331), .B(n330), .C(n535), .Y(n332) );
  NAND2XL U139 ( .A(n101), .B(n31), .Y(n326) );
  NAND2XL U140 ( .A(n98), .B(n103), .Y(n325) );
  NAND2XL U141 ( .A(n87), .B(n15), .Y(n419) );
  NAND2XL U142 ( .A(n15), .B(n92), .Y(n141) );
  NAND2XL U143 ( .A(n104), .B(b[4]), .Y(n510) );
  NAND2XL U144 ( .A(n97), .B(n25), .Y(n416) );
  NAND2XL U145 ( .A(n104), .B(n96), .Y(n514) );
  NAND2XL U146 ( .A(n32), .B(n103), .Y(n513) );
  NAND2XL U147 ( .A(n95), .B(n21), .Y(n420) );
  NAND2XL U148 ( .A(n107), .B(n31), .Y(n454) );
  NAND2XL U149 ( .A(n5), .B(n102), .Y(n319) );
  NAND2XL U150 ( .A(n101), .B(n6), .Y(n290) );
  NAND2XL U151 ( .A(n32), .B(n101), .Y(n493) );
  NAND2XL U152 ( .A(n21), .B(n33), .Y(n246) );
  NAND2XL U153 ( .A(n105), .B(b[4]), .Y(n522) );
  XOR2X1 U154 ( .A(n203), .B(n202), .Y(n204) );
  NAND2XL U155 ( .A(n14), .B(n100), .Y(n85) );
  NAND2XL U156 ( .A(n96), .B(n15), .Y(n449) );
  NAND2XL U157 ( .A(n20), .B(n100), .Y(n298) );
  NAND2XL U158 ( .A(n106), .B(n100), .Y(n195) );
  NAND2XL U159 ( .A(n30), .B(n20), .Y(n194) );
  NAND2XL U160 ( .A(n105), .B(n100), .Y(n468) );
  NAND2XL U161 ( .A(n97), .B(n104), .Y(n320) );
  NAND2XL U162 ( .A(n96), .B(n102), .Y(n494) );
  NAND2XL U163 ( .A(n23), .B(n99), .Y(n481) );
  NAND2XL U164 ( .A(n105), .B(n32), .Y(n337) );
  NAND2XL U165 ( .A(n31), .B(n102), .Y(n339) );
  NAND2XL U166 ( .A(n98), .B(n23), .Y(n440) );
  NAND2XL U167 ( .A(n97), .B(n23), .Y(n396) );
  NAND2XL U168 ( .A(n95), .B(n107), .Y(n404) );
  NAND2XL U169 ( .A(a[5]), .B(n10), .Y(n335) );
  NAND2BXL U170 ( .AN(b[11]), .B(a[12]), .Y(n108) );
  NAND2XL U171 ( .A(n11), .B(n18), .Y(n421) );
  NAND2XL U172 ( .A(n23), .B(n5), .Y(n455) );
  NAND2XL U173 ( .A(n103), .B(n95), .Y(n501) );
  NAND2XL U174 ( .A(n98), .B(n14), .Y(n193) );
  NAND2XL U175 ( .A(n4), .B(n18), .Y(n192) );
  AOI22XL U176 ( .A0(n15), .A1(n410), .B0(n37), .B1(n409), .Y(n412) );
  NAND2XL U177 ( .A(n11), .B(n21), .Y(n414) );
  XNOR2X1 U178 ( .A(n52), .B(n321), .Y(n323) );
  NAND2XL U179 ( .A(n24), .B(n87), .Y(n52) );
  NAND2XL U180 ( .A(n96), .B(n101), .Y(n53) );
  XOR3X2 U181 ( .A(n54), .B(n304), .C(n334), .Y(n305) );
  NAND2XL U182 ( .A(n32), .B(n102), .Y(n54) );
  OAI2BB1XL U183 ( .A0N(n37), .A1N(n188), .B0(n86), .Y(n191) );
  AOI22XL U184 ( .A0(n25), .A1(n507), .B0(n24), .B1(n506), .Y(n509) );
  NAND2XL U185 ( .A(n86), .B(n299), .Y(n302) );
  NAND2BXL U186 ( .AN(n5), .B(n37), .Y(n299) );
  NAND2XL U187 ( .A(n101), .B(b[4]), .Y(n213) );
  NAND2XL U188 ( .A(n97), .B(n20), .Y(n77) );
  NAND2XL U189 ( .A(n17), .B(n96), .Y(n81) );
  NAND2XL U190 ( .A(n12), .B(n102), .Y(n128) );
  NAND2XL U191 ( .A(b[11]), .B(n103), .Y(n131) );
  NAND2XL U192 ( .A(n20), .B(n96), .Y(n83) );
  NAND2XL U193 ( .A(n17), .B(n95), .Y(n84) );
  AOI22XL U194 ( .A0(n24), .A1(n517), .B0(n21), .B1(n516), .Y(n521) );
  NAND2XL U195 ( .A(n101), .B(n12), .Y(n426) );
  NAND2XL U196 ( .A(n96), .B(n24), .Y(n417) );
  NAND2XL U197 ( .A(n33), .B(n15), .Y(n408) );
  AND2X1 U198 ( .A(n36), .B(n100), .Y(n64) );
  NAND2XL U199 ( .A(n106), .B(n30), .Y(n442) );
  NAND2XL U200 ( .A(n107), .B(n4), .Y(n439) );
  INVXL U201 ( .A(n100), .Y(n386) );
  AND2X1 U202 ( .A(n15), .B(n95), .Y(n151) );
  AND2X1 U203 ( .A(n97), .B(n14), .Y(n177) );
  AND2X1 U204 ( .A(n17), .B(n99), .Y(n240) );
  AND2X1 U205 ( .A(n105), .B(n96), .Y(n321) );
  INVXL U206 ( .A(n95), .Y(n170) );
  NAND2XL U207 ( .A(n15), .B(n99), .Y(n55) );
  XNOR2X1 U208 ( .A(n298), .B(n297), .Y(n57) );
  XOR2X1 U209 ( .A(n453), .B(n452), .Y(n461) );
  XOR2X1 U210 ( .A(n451), .B(n450), .Y(n452) );
  NAND2XL U211 ( .A(n97), .B(n18), .Y(n451) );
  NAND2XL U212 ( .A(n5), .B(n103), .Y(n347) );
  NAND2XL U213 ( .A(n101), .B(n33), .Y(n357) );
  NAND2XL U214 ( .A(n25), .B(n10), .Y(n353) );
  NAND2XL U215 ( .A(a[5]), .B(n32), .Y(n354) );
  NAND2XL U216 ( .A(n26), .B(n6), .Y(n355) );
  NAND2XL U217 ( .A(b[4]), .B(n24), .Y(n413) );
  NAND2XL U218 ( .A(n27), .B(n31), .Y(n429) );
  NAND2XL U219 ( .A(n27), .B(n5), .Y(n407) );
  NAND2XL U220 ( .A(b[4]), .B(n102), .Y(n486) );
  NAND2XL U221 ( .A(a[1]), .B(n33), .Y(n431) );
  AND2X1 U222 ( .A(n21), .B(n87), .Y(n402) );
  NAND2XL U223 ( .A(n28), .B(n31), .Y(n406) );
  AND2X1 U224 ( .A(n5), .B(a[0]), .Y(n528) );
  NAND2XL U225 ( .A(n11), .B(n102), .Y(n211) );
  NAND2XL U226 ( .A(n106), .B(n11), .Y(n523) );
  NAND2XL U227 ( .A(n28), .B(b[10]), .Y(n432) );
  NAND2XL U228 ( .A(a[1]), .B(b[10]), .Y(n356) );
  NAND2XL U229 ( .A(n26), .B(n5), .Y(n430) );
  NAND2XL U230 ( .A(n86), .B(n135), .Y(n138) );
  NAND2BXL U231 ( .AN(b[1]), .B(a[11]), .Y(n135) );
  AOI2BB2XL U232 ( .B0(b[0]), .B1(n373), .A0N(n86), .A1N(n366), .Y(n368) );
  INVXL U233 ( .A(b[1]), .Y(n366) );
  XNOR2X1 U234 ( .A(n43), .B(n375), .Y(n288) );
  XOR2X1 U235 ( .A(n61), .B(n381), .Y(n266) );
  XOR3X2 U236 ( .A(n263), .B(n262), .C(n261), .Y(n264) );
  XNOR3X2 U237 ( .A(n180), .B(n43), .C(n179), .Y(n182) );
  XOR3X2 U238 ( .A(n512), .B(n38), .C(n382), .Y(n389) );
  XNOR3X2 U239 ( .A(n43), .B(n505), .C(n216), .Y(n286) );
  XOR2X1 U240 ( .A(n495), .B(n64), .Y(n216) );
  XOR2X1 U241 ( .A(n504), .B(n503), .Y(n505) );
  XOR2X1 U242 ( .A(n494), .B(n493), .Y(n495) );
  XOR3X2 U243 ( .A(n360), .B(n359), .C(n358), .Y(n361) );
  XOR2X1 U244 ( .A(n406), .B(n407), .Y(n359) );
  XNOR3X2 U245 ( .A(n413), .B(n357), .C(n356), .Y(n358) );
  XOR2X1 U246 ( .A(n377), .B(n64), .Y(n360) );
  XNOR3X2 U247 ( .A(n177), .B(n176), .C(n175), .Y(n178) );
  INVX1 U248 ( .A(n382), .Y(n375) );
  XOR2X1 U249 ( .A(n286), .B(n266), .Y(c[6]) );
  XOR2X1 U250 ( .A(n436), .B(n435), .Y(c[12]) );
  XNOR2X1 U251 ( .A(n296), .B(n38), .Y(n61) );
  XOR2X1 U252 ( .A(n527), .B(n526), .Y(n529) );
  XOR2X1 U253 ( .A(n525), .B(n524), .Y(n526) );
  XOR2X1 U254 ( .A(n389), .B(n515), .Y(n527) );
  XOR2X1 U255 ( .A(n523), .B(n522), .Y(n524) );
  XOR2X1 U256 ( .A(n475), .B(n470), .Y(n187) );
  XOR2X1 U257 ( .A(n474), .B(n473), .Y(n475) );
  NOR2X1 U258 ( .A(n384), .B(n519), .Y(n473) );
  XOR3X2 U259 ( .A(n180), .B(n179), .C(n376), .Y(n63) );
  XNOR3X2 U260 ( .A(n63), .B(n215), .C(n214), .Y(c[4]) );
  XOR3X2 U261 ( .A(n352), .B(n528), .C(n529), .Y(c[8]) );
  XNOR2X1 U262 ( .A(n306), .B(n305), .Y(c[7]) );
  XOR3X2 U263 ( .A(n187), .B(n182), .C(n181), .Y(c[3]) );
  XNOR3X2 U264 ( .A(n333), .B(n61), .C(n332), .Y(c[9]) );
  NOR2X1 U265 ( .A(n519), .B(n383), .Y(n508) );
  OAI21XL U266 ( .A0(n33), .A1(n365), .B0(n86), .Y(n127) );
  OAI21XL U267 ( .A0(n18), .A1(n531), .B0(n8), .Y(n534) );
  OAI21XL U268 ( .A0(n21), .A1(n9), .B0(n7), .Y(n533) );
  AOI22X1 U269 ( .A0(n103), .A1(n472), .B0(n104), .B1(n471), .Y(n474) );
  OAI21XL U270 ( .A0(n104), .A1(n366), .B0(n59), .Y(n472) );
  OAI21XL U271 ( .A0(n103), .A1(n9), .B0(n7), .Y(n471) );
  AOI22X1 U272 ( .A0(n15), .A1(n401), .B0(n18), .B1(n400), .Y(n403) );
  OAI21XL U273 ( .A0(n18), .A1(n9), .B0(n58), .Y(n401) );
  INVXL U274 ( .A(n97), .Y(n252) );
  OAI2BB1X1 U275 ( .A0N(n31), .A1N(n317), .B0(n316), .Y(n318) );
  OAI21XL U276 ( .A0(n21), .A1(n366), .B0(n59), .Y(n517) );
  OAI21XL U277 ( .A0(n26), .A1(n366), .B0(n8), .Y(n477) );
  OAI21XL U278 ( .A0(n24), .A1(n366), .B0(n8), .Y(n507) );
  OAI21XL U279 ( .A0(n37), .A1(n366), .B0(n59), .Y(n410) );
  OAI21XL U280 ( .A0(n106), .A1(n9), .B0(n58), .Y(n496) );
  OAI21XL U281 ( .A0(n24), .A1(n9), .B0(n7), .Y(n516) );
  OAI21XL U282 ( .A0(n102), .A1(n532), .B0(n7), .Y(n444) );
  OAI21XL U283 ( .A0(n27), .A1(n532), .B0(n7), .Y(n476) );
  AOI22X1 U284 ( .A0(n26), .A1(n483), .B0(a[5]), .B1(n482), .Y(n484) );
  OAI21XL U285 ( .A0(a[5]), .A1(n366), .B0(n8), .Y(n483) );
  OAI21XL U286 ( .A0(n105), .A1(n9), .B0(n7), .Y(n482) );
  OAI21XL U287 ( .A0(n25), .A1(n9), .B0(n7), .Y(n506) );
  OAI21XL U288 ( .A0(n15), .A1(n9), .B0(n7), .Y(n409) );
  INVX1 U289 ( .A(n87), .Y(n519) );
  OAI2BB1X1 U290 ( .A0N(a[11]), .A1N(n95), .B0(n388), .Y(n372) );
  XNOR3X2 U291 ( .A(n441), .B(n163), .C(n162), .Y(n164) );
  XNOR3X2 U292 ( .A(n151), .B(n150), .C(n149), .Y(n165) );
  NAND2X1 U293 ( .A(n105), .B(n99), .Y(n441) );
  XNOR3X2 U294 ( .A(n395), .B(n134), .C(n133), .Y(n143) );
  XNOR3X2 U295 ( .A(n141), .B(n140), .C(n139), .Y(n142) );
  XNOR2X1 U296 ( .A(n481), .B(n480), .Y(n205) );
  XOR2X1 U297 ( .A(n247), .B(n246), .Y(n248) );
  XNOR3X2 U298 ( .A(n240), .B(n239), .C(n221), .Y(n249) );
  NOR2X1 U299 ( .A(n386), .B(n462), .Y(n463) );
  XOR2X1 U300 ( .A(n461), .B(n460), .Y(n464) );
  INVX1 U301 ( .A(n104), .Y(n462) );
  AOI21XL U302 ( .A0(n37), .A1(n170), .B0(n370), .Y(n174) );
  NAND2X1 U303 ( .A(n107), .B(n100), .Y(n262) );
  NOR2BX1 U304 ( .AN(a[12]), .B(n87), .Y(n136) );
  OAI21XL U305 ( .A0(n146), .A1(n373), .B0(n87), .Y(n147) );
  NAND2X1 U306 ( .A(n105), .B(n33), .Y(n456) );
  NAND2X1 U307 ( .A(n23), .B(b[11]), .Y(n250) );
  XOR2X1 U308 ( .A(n502), .B(n501), .Y(n503) );
  XNOR2X1 U309 ( .A(n193), .B(n192), .Y(n203) );
  XOR3X2 U310 ( .A(n378), .B(n380), .C(n381), .Y(n490) );
  XOR2X1 U311 ( .A(n375), .B(n38), .Y(n380) );
  XOR2X1 U312 ( .A(n291), .B(n290), .Y(n304) );
  NAND2X1 U313 ( .A(n10), .B(n103), .Y(n291) );
  XOR2X1 U314 ( .A(n447), .B(n446), .Y(n465) );
  NOR2X1 U315 ( .A(n385), .B(n519), .Y(n446) );
  AOI22X1 U316 ( .A0(n102), .A1(n445), .B0(n28), .B1(n444), .Y(n447) );
  OAI21XL U317 ( .A0(n28), .A1(n366), .B0(n8), .Y(n445) );
  XOR2X1 U318 ( .A(n168), .B(n167), .Y(n176) );
  XOR2X1 U319 ( .A(n153), .B(n152), .Y(n163) );
  XOR2X1 U320 ( .A(n397), .B(n398), .Y(n134) );
  NAND2BX1 U321 ( .AN(n97), .B(a[11]), .Y(n254) );
  XOR2X1 U322 ( .A(n195), .B(n194), .Y(n202) );
  XOR2X1 U323 ( .A(n459), .B(n458), .Y(n460) );
  XOR2X1 U324 ( .A(n455), .B(n454), .Y(n459) );
  XOR2X1 U325 ( .A(n457), .B(n456), .Y(n458) );
  XOR2X1 U326 ( .A(n423), .B(n422), .Y(n424) );
  XOR2X1 U327 ( .A(n421), .B(n420), .Y(n422) );
  XOR2X1 U328 ( .A(n369), .B(n419), .Y(n423) );
  XNOR3X2 U329 ( .A(n509), .B(n289), .C(n288), .Y(n306) );
  XOR3X2 U330 ( .A(n510), .B(n511), .C(n508), .Y(n289) );
  XNOR3X2 U331 ( .A(n412), .B(n352), .C(n351), .Y(n363) );
  XNOR2X1 U332 ( .A(n411), .B(n414), .Y(n351) );
  NAND2X1 U333 ( .A(n4), .B(n14), .Y(n251) );
  NAND2X1 U334 ( .A(n106), .B(n99), .Y(n457) );
  XNOR3X2 U335 ( .A(n324), .B(n323), .C(n538), .Y(n333) );
  XOR2X1 U336 ( .A(n320), .B(n319), .Y(n324) );
  OAI2BB1X1 U337 ( .A0N(n31), .A1N(n302), .B0(n301), .Y(n303) );
  OAI21XL U338 ( .A0(n300), .A1(n373), .B0(n5), .Y(n301) );
  XNOR3X2 U339 ( .A(n77), .B(n81), .C(n440), .Y(n149) );
  XNOR3X2 U340 ( .A(n83), .B(n84), .C(n396), .Y(n139) );
  XOR3X2 U341 ( .A(n536), .B(n537), .C(n327), .Y(n331) );
  XNOR3X2 U342 ( .A(n479), .B(n213), .C(n212), .Y(n214) );
  XOR2X1 U343 ( .A(n211), .B(n478), .Y(n212) );
  AOI22X1 U344 ( .A0(n27), .A1(n477), .B0(n26), .B1(n476), .Y(n479) );
  XNOR3X2 U345 ( .A(n132), .B(n131), .C(n128), .Y(n133) );
  NAND2X1 U346 ( .A(n30), .B(n17), .Y(n263) );
  NAND2X1 U347 ( .A(n107), .B(n99), .Y(n466) );
  XOR2X2 U348 ( .A(n111), .B(n85), .Y(n144) );
  OAI2BB1X1 U349 ( .A0N(n5), .A1N(n220), .B0(n219), .Y(n221) );
  OAI21XL U350 ( .A0(n217), .A1(n373), .B0(n98), .Y(n219) );
  XNOR3X2 U351 ( .A(n399), .B(n350), .C(n179), .Y(c[0]) );
  XOR2X1 U352 ( .A(n500), .B(n499), .Y(n504) );
  NOR2X1 U353 ( .A(n519), .B(n498), .Y(n499) );
  AOI22X1 U354 ( .A0(n106), .A1(n497), .B0(n107), .B1(n496), .Y(n500) );
  INVX1 U355 ( .A(n105), .Y(n498) );
  XOR2X1 U356 ( .A(n521), .B(n520), .Y(n525) );
  NOR2X1 U357 ( .A(n519), .B(n518), .Y(n520) );
  INVX1 U358 ( .A(n107), .Y(n518) );
  XOR2X1 U359 ( .A(n428), .B(n427), .Y(n436) );
  XNOR2X1 U360 ( .A(n426), .B(n538), .Y(n427) );
  XOR2X1 U361 ( .A(n425), .B(n424), .Y(n428) );
  XOR2X1 U362 ( .A(n449), .B(n448), .Y(n453) );
  XOR2X1 U363 ( .A(n394), .B(n418), .Y(n425) );
  XOR2X1 U364 ( .A(n417), .B(n416), .Y(n418) );
  XOR2X1 U365 ( .A(n364), .B(n415), .Y(n394) );
  XOR2X1 U366 ( .A(n489), .B(n488), .Y(n491) );
  XOR2X1 U367 ( .A(n487), .B(n486), .Y(n488) );
  XOR2X1 U368 ( .A(n485), .B(n484), .Y(n489) );
  NAND2X1 U369 ( .A(n28), .B(n11), .Y(n487) );
  NAND2BX1 U370 ( .AN(n98), .B(n36), .Y(n253) );
  XNOR2X1 U371 ( .A(n442), .B(n439), .Y(n162) );
  XOR2X1 U372 ( .A(n468), .B(n469), .Y(n166) );
  AOI22X1 U373 ( .A0(a[0]), .A1(n438), .B0(a[1]), .B1(n437), .Y(n443) );
  OAI21XL U374 ( .A0(a[1]), .A1(n531), .B0(n8), .Y(n438) );
  OAI21XL U375 ( .A0(n101), .A1(n9), .B0(n7), .Y(n437) );
  NOR2X1 U376 ( .A(n519), .B(n530), .Y(n478) );
  INVX1 U377 ( .A(n103), .Y(n530) );
  NOR2X1 U378 ( .A(n385), .B(n9), .Y(n399) );
  XOR2X1 U379 ( .A(n514), .B(n513), .Y(n515) );
  XOR2X1 U380 ( .A(n434), .B(n433), .Y(n435) );
  XOR2X1 U381 ( .A(n430), .B(n429), .Y(n434) );
  XOR2X1 U382 ( .A(n432), .B(n431), .Y(n433) );
  NAND2X1 U383 ( .A(n27), .B(n87), .Y(n485) );
  XOR3X2 U384 ( .A(n339), .B(n338), .C(n337), .Y(n346) );
  NAND2X1 U385 ( .A(n101), .B(b[10]), .Y(n338) );
  XNOR3X2 U386 ( .A(n355), .B(n354), .C(n353), .Y(n362) );
  INVX1 U387 ( .A(n101), .Y(n385) );
  XOR2X1 U388 ( .A(n326), .B(n325), .Y(n327) );
  XOR2X1 U389 ( .A(n405), .B(n404), .Y(n348) );
  INVX1 U390 ( .A(n102), .Y(n384) );
  INVX1 U391 ( .A(n106), .Y(n383) );
  OAI2BB1X1 U392 ( .A0N(n87), .A1N(n138), .B0(n137), .Y(n140) );
  OAI21XL U393 ( .A0(n136), .A1(n373), .B0(b[1]), .Y(n137) );
  BUFX3 U394 ( .A(a[3]), .Y(n104) );
  BUFX3 U395 ( .A(a[6]), .Y(n107) );
  BUFX3 U396 ( .A(a[2]), .Y(n103) );
  BUFX3 U397 ( .A(a[4]), .Y(n105) );
  BUFX3 U398 ( .A(a[5]), .Y(n106) );
  BUFX3 U399 ( .A(a[1]), .Y(n102) );
  BUFX3 U400 ( .A(b[12]), .Y(n100) );
  BUFX3 U401 ( .A(b[7]), .Y(n98) );
  INVX1 U402 ( .A(b[0]), .Y(n532) );
  INVX1 U403 ( .A(b[1]), .Y(n531) );
  BUFX3 U404 ( .A(b[2]), .Y(n87) );
  BUFX3 U405 ( .A(a[0]), .Y(n101) );
  OAI21XL U406 ( .A0(n100), .A1(n34), .B0(n311), .Y(n122) );
  XOR2X1 U407 ( .A(n144), .B(n377), .Y(n350) );
endmodule


module multiplier_11 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n47, n49, n50, n51, n52,
         n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n74, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n92,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n122, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n202,
         n203, n204, n205, n210, n211, n212, n213, n214, n215, n216, n217,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n230,
         n233, n234, n235, n236, n237, n238, n239, n240, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n259, n260, n261, n262, n263,
         n264, n265, n266, n278, n286, n288, n289, n290, n291, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n311, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n343, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503;

  CLKINVX3 U1 ( .A(n316), .Y(n381) );
  OAI21XL U2 ( .A0(n381), .A1(n143), .B0(n86), .Y(n144) );
  OAI211X1 U3 ( .A0(n377), .A1(n60), .B0(n383), .C0(n382), .Y(n384) );
  XOR2X1 U4 ( .A(n385), .B(n5), .Y(n362) );
  OAI2BB1X1 U5 ( .A0N(n99), .A1N(n107), .B0(n106), .Y(n109) );
  NOR2X1 U6 ( .A(n188), .B(n189), .Y(n1) );
  INVXL U7 ( .A(n1), .Y(n190) );
  OAI21XL U8 ( .A0(n2), .A1(n322), .B0(n323), .Y(n324) );
  INVX1 U9 ( .A(n321), .Y(n2) );
  NOR2X1 U10 ( .A(n490), .B(n24), .Y(n455) );
  NOR2XL U11 ( .A(n490), .B(n14), .Y(n408) );
  OAI21XL U12 ( .A0(n3), .A1(n98), .B0(n316), .Y(n318) );
  INVX1 U13 ( .A(n39), .Y(n3) );
  OR2X2 U14 ( .A(n189), .B(n181), .Y(n192) );
  AND2X2 U15 ( .A(n86), .B(n104), .Y(n491) );
  NOR2X1 U16 ( .A(n24), .B(n320), .Y(n84) );
  XNOR2X1 U17 ( .A(n221), .B(n439), .Y(c[1]) );
  NAND3X1 U18 ( .A(n189), .B(n181), .C(n188), .Y(n191) );
  AOI211XL U19 ( .A0(n318), .A1(n34), .B0(n323), .C0(n32), .Y(n4) );
  INVX1 U20 ( .A(n4), .Y(n326) );
  OAI2BB1X1 U21 ( .A0N(a[11]), .A1N(n320), .B0(n85), .Y(n107) );
  XOR2X2 U22 ( .A(n109), .B(n108), .Y(n375) );
  OAI21XL U23 ( .A0(n105), .A1(n381), .B0(n98), .Y(n106) );
  XOR2X2 U24 ( .A(n263), .B(n66), .Y(n278) );
  XOR2X2 U25 ( .A(n195), .B(n194), .Y(n263) );
  XNOR3X2 U26 ( .A(n52), .B(n53), .C(n301), .Y(n5) );
  AND2X2 U27 ( .A(n101), .B(n34), .Y(n6) );
  XNOR3X2 U28 ( .A(n238), .B(n237), .C(n236), .Y(n7) );
  NAND2X1 U29 ( .A(b[1]), .B(n497), .Y(n8) );
  INVX1 U30 ( .A(b[12]), .Y(n9) );
  INVX1 U31 ( .A(n9), .Y(n10) );
  CLKINVX2 U32 ( .A(n9), .Y(n11) );
  INVX1 U33 ( .A(n388), .Y(n12) );
  INVX1 U34 ( .A(n214), .Y(n13) );
  INVX1 U35 ( .A(a[9]), .Y(n14) );
  INVX1 U36 ( .A(n14), .Y(n15) );
  INVX1 U37 ( .A(n14), .Y(n16) );
  INVX1 U38 ( .A(a[8]), .Y(n17) );
  INVX1 U39 ( .A(n17), .Y(n18) );
  INVX1 U40 ( .A(a[7]), .Y(n19) );
  INVXL U41 ( .A(n19), .Y(n20) );
  INVX1 U42 ( .A(a[3]), .Y(n21) );
  INVXL U43 ( .A(n21), .Y(n22) );
  INVX1 U44 ( .A(n495), .Y(n23) );
  INVX1 U45 ( .A(a[1]), .Y(n24) );
  INVX1 U46 ( .A(n24), .Y(n25) );
  INVX1 U47 ( .A(n110), .Y(n26) );
  INVX1 U48 ( .A(b[8]), .Y(n27) );
  INVX1 U49 ( .A(n27), .Y(n28) );
  INVX1 U50 ( .A(n225), .Y(n29) );
  INVX1 U51 ( .A(n164), .Y(n30) );
  INVX1 U52 ( .A(n389), .Y(n31) );
  INVX1 U53 ( .A(n320), .Y(n32) );
  INVX1 U54 ( .A(b[9]), .Y(n33) );
  INVX1 U55 ( .A(n33), .Y(n34) );
  XOR2X2 U56 ( .A(n264), .B(n174), .Y(n202) );
  NAND2BX1 U57 ( .AN(a[12]), .B(a[11]), .Y(n380) );
  BUFX3 U58 ( .A(n380), .Y(n85) );
  NAND2X1 U59 ( .A(b[0]), .B(n496), .Y(n35) );
  NAND2X1 U60 ( .A(b[0]), .B(n496), .Y(n61) );
  INVX1 U61 ( .A(a[10]), .Y(n36) );
  INVX1 U62 ( .A(n36), .Y(n37) );
  INVXL U63 ( .A(n36), .Y(n38) );
  AND2X1 U64 ( .A(n37), .B(n10), .Y(n108) );
  BUFX3 U65 ( .A(a[12]), .Y(n39) );
  INVX1 U66 ( .A(n377), .Y(n47) );
  INVX1 U67 ( .A(b[0]), .Y(n49) );
  NAND2XL U68 ( .A(n15), .B(n10), .Y(n315) );
  NAND2X1 U69 ( .A(n37), .B(n99), .Y(n314) );
  XNOR3X2 U70 ( .A(n173), .B(n50), .C(n51), .Y(n264) );
  XNOR3X2 U71 ( .A(n155), .B(n446), .C(n79), .Y(n50) );
  XNOR3X2 U72 ( .A(n170), .B(n169), .C(n168), .Y(n51) );
  INVXL U73 ( .A(n375), .Y(n141) );
  NOR2XL U74 ( .A(n59), .B(n320), .Y(n322) );
  INVXL U75 ( .A(n323), .Y(n319) );
  XOR2X1 U76 ( .A(n74), .B(n447), .Y(c[2]) );
  INVXL U77 ( .A(n99), .Y(n110) );
  OAI2BB1XL U78 ( .A0N(n47), .A1N(n110), .B0(n85), .Y(n126) );
  AOI22XL U79 ( .A0(n23), .A1(n454), .B0(n22), .B1(n453), .Y(n456) );
  AOI22XL U80 ( .A0(n18), .A1(n499), .B0(n16), .B1(n498), .Y(n501) );
  NAND2XL U81 ( .A(n97), .B(n104), .Y(n395) );
  AOI22XL U82 ( .A0(n38), .A1(n401), .B0(n16), .B1(n400), .Y(n402) );
  NAND2XL U83 ( .A(n30), .B(a[6]), .Y(n403) );
  NAND2XL U84 ( .A(n28), .B(n38), .Y(n234) );
  NAND2XL U85 ( .A(b[9]), .B(n38), .Y(n253) );
  NAND2XL U86 ( .A(n103), .B(n98), .Y(n446) );
  NAND2BXL U87 ( .AN(n97), .B(n47), .Y(n248) );
  NAND2XL U88 ( .A(n85), .B(n248), .Y(n251) );
  NAND2BXL U89 ( .AN(n86), .B(a[11]), .Y(n142) );
  NAND2XL U90 ( .A(n85), .B(n142), .Y(n145) );
  NAND2BXL U91 ( .AN(n96), .B(n39), .Y(n215) );
  NAND2XL U92 ( .A(n38), .B(n98), .Y(n52) );
  XNOR2X1 U93 ( .A(n296), .B(n291), .Y(n53) );
  NAND2XL U94 ( .A(n10), .B(n101), .Y(n150) );
  NAND2XL U95 ( .A(a[3]), .B(n99), .Y(n149) );
  NAND2XL U96 ( .A(n102), .B(b[9]), .Y(n397) );
  NAND2XL U97 ( .A(n103), .B(b[8]), .Y(n398) );
  NOR2X1 U98 ( .A(n230), .B(n228), .Y(n237) );
  AOI21XL U99 ( .A0(n85), .A1(n227), .B0(n388), .Y(n228) );
  NAND2XL U100 ( .A(a[7]), .B(n34), .Y(n449) );
  NAND2XL U101 ( .A(n39), .B(n11), .Y(n366) );
  NAND2XL U102 ( .A(n86), .B(n38), .Y(n416) );
  NAND2BXL U103 ( .AN(b[8]), .B(n47), .Y(n297) );
  NAND2XL U104 ( .A(n85), .B(n297), .Y(n300) );
  NAND2XL U105 ( .A(n20), .B(n26), .Y(n233) );
  XOR2X1 U106 ( .A(n154), .B(n153), .Y(n175) );
  NAND2XL U107 ( .A(n102), .B(n98), .Y(n437) );
  AOI22XL U108 ( .A0(n20), .A1(n489), .B0(n18), .B1(n488), .Y(n492) );
  NAND2XL U109 ( .A(n29), .B(n23), .Y(n78) );
  NAND2XL U110 ( .A(a[4]), .B(n13), .Y(n334) );
  NAND2XL U111 ( .A(n87), .B(n20), .Y(n404) );
  NAND2XL U112 ( .A(n104), .B(n98), .Y(n448) );
  NAND2XL U113 ( .A(a[3]), .B(n92), .Y(n486) );
  NAND2XL U114 ( .A(n96), .B(n37), .Y(n177) );
  NAND2XL U115 ( .A(b[8]), .B(a[8]), .Y(n178) );
  NAND2XL U116 ( .A(n97), .B(n15), .Y(n179) );
  NAND2XL U117 ( .A(b[9]), .B(n16), .Y(n235) );
  NAND2XL U118 ( .A(n34), .B(n318), .Y(n321) );
  NAND2XL U119 ( .A(n30), .B(a[1]), .Y(n467) );
  INVXL U120 ( .A(n97), .Y(n388) );
  NAND2XL U121 ( .A(n103), .B(n11), .Y(n212) );
  NAND2XL U122 ( .A(n96), .B(n104), .Y(n413) );
  NAND2XL U123 ( .A(n104), .B(b[8]), .Y(n435) );
  NAND2XL U124 ( .A(n103), .B(b[9]), .Y(n438) );
  NAND2XL U125 ( .A(a[7]), .B(n32), .Y(n462) );
  NAND2XL U126 ( .A(n101), .B(n92), .Y(n477) );
  NAND2XL U127 ( .A(n15), .B(n99), .Y(n291) );
  NAND2XL U128 ( .A(n18), .B(n26), .Y(n259) );
  NAND2XL U129 ( .A(n104), .B(n11), .Y(n223) );
  NAND2XL U130 ( .A(a[7]), .B(b[8]), .Y(n445) );
  NOR2BXL U131 ( .AN(n39), .B(n11), .Y(n111) );
  NAND2XL U132 ( .A(n31), .B(a[6]), .Y(n503) );
  NAND2XL U133 ( .A(n97), .B(n38), .Y(n213) );
  NAND2XL U134 ( .A(n18), .B(n98), .Y(n224) );
  NAND2XL U135 ( .A(n101), .B(n31), .Y(n468) );
  NAND2XL U136 ( .A(n104), .B(n99), .Y(n461) );
  NAND2XL U137 ( .A(a[8]), .B(n10), .Y(n296) );
  AND2X1 U138 ( .A(n87), .B(a[1]), .Y(n205) );
  INVXL U139 ( .A(n103), .Y(n386) );
  XNOR3X2 U140 ( .A(n54), .B(n55), .C(n219), .Y(n220) );
  NAND2XL U141 ( .A(n34), .B(n18), .Y(n54) );
  NAND2XL U142 ( .A(n28), .B(n16), .Y(n55) );
  NAND2XL U143 ( .A(n97), .B(a[7]), .Y(n436) );
  NAND2XL U144 ( .A(n96), .B(a[7]), .Y(n396) );
  NAND2BXL U145 ( .AN(n96), .B(a[11]), .Y(n227) );
  NAND2XL U146 ( .A(n97), .B(n22), .Y(n355) );
  NAND2XL U147 ( .A(n103), .B(n95), .Y(n354) );
  NAND2XL U148 ( .A(n87), .B(n16), .Y(n418) );
  NAND2XL U149 ( .A(n92), .B(n18), .Y(n417) );
  NAND2XL U150 ( .A(n95), .B(a[1]), .Y(n470) );
  NAND2XL U151 ( .A(n96), .B(n100), .Y(n469) );
  AOI22XL U152 ( .A0(n38), .A1(n407), .B0(n47), .B1(n406), .Y(n409) );
  NAND2XL U153 ( .A(n31), .B(n18), .Y(n411) );
  OAI2BB1XL U154 ( .A0N(n47), .A1N(n214), .B0(n85), .Y(n217) );
  XOR3X2 U155 ( .A(n57), .B(n302), .C(n360), .Y(n303) );
  NAND2XL U156 ( .A(n29), .B(n25), .Y(n57) );
  NAND2XL U157 ( .A(n100), .B(n11), .Y(n423) );
  AOI22XL U158 ( .A0(a[6]), .A1(n483), .B0(n20), .B1(n482), .Y(n485) );
  NAND2XL U159 ( .A(n102), .B(n31), .Y(n487) );
  INVXL U160 ( .A(n87), .Y(n389) );
  XOR3X2 U161 ( .A(n58), .B(n353), .C(n352), .Y(n357) );
  NAND2XL U162 ( .A(n18), .B(n86), .Y(n58) );
  NAND2XL U163 ( .A(n11), .B(a[1]), .Y(n134) );
  NAND2XL U164 ( .A(n99), .B(n101), .Y(n135) );
  NAND2XL U165 ( .A(n98), .B(a[3]), .Y(n136) );
  NOR2BXL U166 ( .AN(a[11]), .B(n92), .Y(n187) );
  NAND2XL U167 ( .A(n96), .B(a[8]), .Y(n82) );
  NAND2XL U168 ( .A(n15), .B(n95), .Y(n83) );
  NAND2XL U169 ( .A(a[8]), .B(n95), .Y(n80) );
  NAND2XL U170 ( .A(n16), .B(n92), .Y(n81) );
  NAND2XL U171 ( .A(n28), .B(n25), .Y(n346) );
  NAND2XL U172 ( .A(a[3]), .B(n87), .Y(n478) );
  NAND2XL U173 ( .A(n95), .B(n20), .Y(n414) );
  XOR2X1 U174 ( .A(n262), .B(n261), .Y(n290) );
  NAND2XL U175 ( .A(n20), .B(n11), .Y(n260) );
  AOI22XL U176 ( .A0(n22), .A1(n458), .B0(n102), .B1(n457), .Y(n460) );
  NAND2XL U177 ( .A(a[5]), .B(n31), .Y(n494) );
  NAND2XL U178 ( .A(n102), .B(n11), .Y(n450) );
  NAND2XL U179 ( .A(n103), .B(n99), .Y(n451) );
  NAND2XL U180 ( .A(n100), .B(n26), .Y(n367) );
  INVXL U181 ( .A(n95), .Y(n214) );
  AND2X1 U182 ( .A(n102), .B(n99), .Y(n79) );
  AND2X1 U183 ( .A(n37), .B(n92), .Y(n148) );
  AND2X1 U184 ( .A(n38), .B(n87), .Y(n133) );
  AND2X1 U185 ( .A(n16), .B(n98), .Y(n254) );
  AND2X1 U186 ( .A(n100), .B(n92), .Y(n210) );
  AND2X1 U187 ( .A(n100), .B(n28), .Y(n327) );
  AND2X1 U188 ( .A(n20), .B(n86), .Y(n500) );
  INVXL U189 ( .A(a[11]), .Y(n377) );
  AND2X1 U190 ( .A(n85), .B(n317), .Y(n59) );
  NAND2XL U191 ( .A(n12), .B(n101), .Y(n338) );
  NAND2XL U192 ( .A(n102), .B(n30), .Y(n493) );
  NAND2XL U193 ( .A(n29), .B(n22), .Y(n337) );
  NAND2XL U194 ( .A(a[6]), .B(n13), .Y(n363) );
  NAND2XL U195 ( .A(a[5]), .B(n29), .Y(n364) );
  NAND2XL U196 ( .A(a[4]), .B(n12), .Y(n365) );
  NAND2XL U197 ( .A(n30), .B(n20), .Y(n410) );
  NAND2XL U198 ( .A(n100), .B(n34), .Y(n339) );
  NAND2XL U199 ( .A(n22), .B(n28), .Y(n405) );
  NAND2XL U200 ( .A(n30), .B(n103), .Y(n502) );
  NAND2XL U201 ( .A(a[4]), .B(n29), .Y(n350) );
  NAND2XL U202 ( .A(n100), .B(n12), .Y(n288) );
  NAND2XL U203 ( .A(n22), .B(n86), .Y(n466) );
  NAND2XL U204 ( .A(n28), .B(n101), .Y(n351) );
  NAND2XL U205 ( .A(a[0]), .B(n13), .Y(n239) );
  NAND2XL U206 ( .A(n13), .B(n22), .Y(n306) );
  NAND2XL U207 ( .A(n12), .B(n25), .Y(n305) );
  NAND2XL U208 ( .A(n23), .B(n32), .Y(n428) );
  NAND2XL U209 ( .A(n25), .B(n26), .Y(n427) );
  NAND2XL U210 ( .A(a[4]), .B(n28), .Y(n426) );
  NAND2XL U211 ( .A(n22), .B(n34), .Y(n425) );
  NAND2BXL U212 ( .AN(b[1]), .B(n47), .Y(n127) );
  NAND2XL U213 ( .A(n85), .B(n127), .Y(n130) );
  INVXL U214 ( .A(b[1]), .Y(n378) );
  NAND2X1 U215 ( .A(b[1]), .B(n497), .Y(n60) );
  XNOR2X1 U216 ( .A(n141), .B(n174), .Y(n359) );
  XNOR2X1 U217 ( .A(n66), .B(n7), .Y(n311) );
  XOR2X1 U218 ( .A(n141), .B(n376), .Y(n62) );
  XOR3X2 U219 ( .A(n360), .B(n359), .C(n358), .Y(c[10]) );
  NAND3X1 U220 ( .A(n326), .B(n325), .C(n324), .Y(n385) );
  NAND3X1 U221 ( .A(n59), .B(n319), .C(n321), .Y(n325) );
  XOR2X1 U222 ( .A(n444), .B(n445), .Y(n173) );
  XNOR3X2 U223 ( .A(n62), .B(n175), .C(n196), .Y(n221) );
  XNOR3X2 U224 ( .A(n333), .B(n332), .C(n331), .Y(c[8]) );
  XOR3X2 U225 ( .A(n202), .B(n263), .C(n196), .Y(n203) );
  XNOR3X2 U226 ( .A(n311), .B(n74), .C(n247), .Y(c[5]) );
  XNOR3X2 U227 ( .A(n465), .B(n246), .C(n240), .Y(n247) );
  XOR2X1 U228 ( .A(n239), .B(n466), .Y(n240) );
  XNOR2X1 U229 ( .A(n468), .B(n467), .Y(n246) );
  INVX1 U230 ( .A(n366), .Y(n376) );
  NOR2X1 U231 ( .A(n386), .B(n388), .Y(n412) );
  XOR3X2 U232 ( .A(n63), .B(n64), .C(n65), .Y(n358) );
  XNOR3X2 U233 ( .A(n404), .B(n403), .C(n402), .Y(n63) );
  XOR2X1 U234 ( .A(n351), .B(n350), .Y(n64) );
  XNOR2X1 U235 ( .A(n357), .B(n356), .Y(n65) );
  INVX1 U236 ( .A(n369), .Y(n174) );
  XOR2X1 U237 ( .A(n224), .B(n223), .Y(n238) );
  XOR3X2 U238 ( .A(n235), .B(n234), .C(n233), .Y(n236) );
  XNOR3X2 U239 ( .A(n376), .B(n264), .C(n263), .Y(n265) );
  XOR3X2 U240 ( .A(n67), .B(n68), .C(n220), .Y(n66) );
  XNOR2X1 U241 ( .A(n213), .B(n212), .Y(n67) );
  XOR2X1 U242 ( .A(n461), .B(n462), .Y(n68) );
  XNOR3X2 U243 ( .A(n77), .B(n266), .C(n265), .Y(c[6]) );
  XOR2X1 U244 ( .A(n481), .B(n471), .Y(n266) );
  XOR2X1 U245 ( .A(n432), .B(n431), .Y(c[12]) );
  XOR2X1 U246 ( .A(n430), .B(n429), .Y(n431) );
  XOR2X1 U247 ( .A(n202), .B(n175), .Y(n74) );
  XOR2X1 U248 ( .A(n371), .B(n370), .Y(n372) );
  XNOR3X2 U249 ( .A(n405), .B(n6), .C(n368), .Y(n371) );
  XOR3X2 U250 ( .A(n410), .B(n369), .C(n84), .Y(n370) );
  INVX1 U251 ( .A(n380), .Y(n182) );
  XNOR2X1 U252 ( .A(n290), .B(n7), .Y(n77) );
  XOR2XL U253 ( .A(n290), .B(n5), .Y(n360) );
  XOR2X1 U254 ( .A(n304), .B(n303), .Y(c[7]) );
  XOR2X1 U255 ( .A(n204), .B(n203), .Y(c[3]) );
  XNOR3X2 U256 ( .A(n77), .B(n349), .C(n348), .Y(c[9]) );
  XOR3X2 U257 ( .A(n374), .B(n373), .C(n372), .Y(c[11]) );
  NOR2XL U258 ( .A(n490), .B(n386), .Y(n484) );
  OAI21XL U259 ( .A0(n16), .A1(n378), .B0(n60), .Y(n499) );
  OAI21XL U260 ( .A0(n18), .A1(n497), .B0(n35), .Y(n498) );
  OAI21XL U261 ( .A0(n22), .A1(n496), .B0(n60), .Y(n454) );
  OAI21XL U262 ( .A0(n101), .A1(n49), .B0(n35), .Y(n453) );
  AOI22X1 U263 ( .A0(n103), .A1(n473), .B0(n104), .B1(n472), .Y(n476) );
  OAI21XL U264 ( .A0(n104), .A1(n378), .B0(n8), .Y(n473) );
  OAI21XL U265 ( .A0(n103), .A1(n497), .B0(n61), .Y(n472) );
  OAI21XL U266 ( .A0(n38), .A1(n378), .B0(n8), .Y(n400) );
  OAI21XL U267 ( .A0(n16), .A1(n49), .B0(n35), .Y(n401) );
  OAI2BB1X1 U268 ( .A0N(n11), .A1N(n126), .B0(n122), .Y(n369) );
  INVXL U269 ( .A(n96), .Y(n225) );
  XNOR3X2 U270 ( .A(n448), .B(n449), .C(n193), .Y(n194) );
  NAND3X1 U271 ( .A(n192), .B(n191), .C(n190), .Y(n195) );
  OAI21XL U272 ( .A0(n25), .A1(n49), .B0(n35), .Y(n440) );
  OAI21XL U273 ( .A0(n22), .A1(n49), .B0(n35), .Y(n457) );
  OAI21XL U274 ( .A0(n20), .A1(n49), .B0(n35), .Y(n488) );
  AOI22X1 U275 ( .A0(a[4]), .A1(n464), .B0(a[5]), .B1(n463), .Y(n465) );
  OAI21XL U276 ( .A0(a[5]), .A1(n378), .B0(n8), .Y(n464) );
  OAI21XL U277 ( .A0(n102), .A1(n49), .B0(n35), .Y(n463) );
  OAI21XL U278 ( .A0(a[6]), .A1(n49), .B0(n35), .Y(n482) );
  OAI21XL U279 ( .A0(n38), .A1(n49), .B0(n35), .Y(n406) );
  OAI21XL U280 ( .A0(n102), .A1(n496), .B0(n60), .Y(n458) );
  OAI21XL U281 ( .A0(n18), .A1(n378), .B0(n8), .Y(n489) );
  OAI21XL U282 ( .A0(n47), .A1(n496), .B0(n60), .Y(n407) );
  XNOR3X2 U283 ( .A(n437), .B(n152), .C(n151), .Y(n153) );
  XNOR3X2 U284 ( .A(n148), .B(n147), .C(n146), .Y(n154) );
  NOR2X1 U285 ( .A(n490), .B(n474), .Y(n475) );
  INVX1 U286 ( .A(n102), .Y(n474) );
  INVX1 U287 ( .A(n86), .Y(n490) );
  OAI2BB1X1 U288 ( .A0N(n87), .A1N(n145), .B0(n144), .Y(n147) );
  XOR2X1 U289 ( .A(n260), .B(n259), .Y(n261) );
  XNOR3X2 U290 ( .A(n254), .B(n253), .C(n252), .Y(n262) );
  NOR2BX1 U291 ( .AN(a[12]), .B(n99), .Y(n105) );
  NOR2BX1 U292 ( .AN(a[11]), .B(n87), .Y(n165) );
  XNOR2X1 U293 ( .A(n315), .B(n314), .Y(n323) );
  XOR2X1 U294 ( .A(n140), .B(n139), .Y(n196) );
  XNOR3X2 U295 ( .A(n395), .B(n138), .C(n137), .Y(n139) );
  XNOR3X2 U296 ( .A(n133), .B(n132), .C(n131), .Y(n140) );
  XNOR3X2 U297 ( .A(n375), .B(n336), .C(n335), .Y(n349) );
  XOR2X1 U298 ( .A(n334), .B(n502), .Y(n335) );
  XNOR2X1 U299 ( .A(n503), .B(n500), .Y(n336) );
  NOR2BX1 U300 ( .AN(a[12]), .B(n95), .Y(n180) );
  XNOR3X2 U301 ( .A(n78), .B(n492), .C(n311), .Y(n332) );
  XNOR3X2 U302 ( .A(n399), .B(n359), .C(n196), .Y(c[0]) );
  XOR2X1 U303 ( .A(n289), .B(n288), .Y(n302) );
  NAND2X1 U304 ( .A(n95), .B(n101), .Y(n289) );
  XNOR3X2 U305 ( .A(n222), .B(n278), .C(n221), .Y(c[4]) );
  XOR2X1 U306 ( .A(n460), .B(n211), .Y(n222) );
  XOR3X2 U307 ( .A(n210), .B(n205), .C(n459), .Y(n211) );
  OAI2BB1X1 U308 ( .A0N(n34), .A1N(n300), .B0(n299), .Y(n301) );
  XOR2X1 U309 ( .A(n163), .B(n162), .Y(n169) );
  NAND2X1 U310 ( .A(n97), .B(a[8]), .Y(n163) );
  NAND2X1 U311 ( .A(n96), .B(n15), .Y(n162) );
  XOR2X1 U312 ( .A(n150), .B(n149), .Y(n152) );
  XOR2X1 U313 ( .A(n397), .B(n398), .Y(n138) );
  XOR3X2 U314 ( .A(n423), .B(n424), .C(n385), .Y(n432) );
  XOR2X1 U315 ( .A(n422), .B(n421), .Y(n424) );
  XOR2X1 U316 ( .A(n420), .B(n419), .Y(n421) );
  XNOR3X2 U317 ( .A(n485), .B(n286), .C(n278), .Y(n304) );
  XOR3X2 U318 ( .A(n486), .B(n487), .C(n484), .Y(n286) );
  XNOR3X2 U319 ( .A(n62), .B(n452), .C(n176), .Y(n204) );
  NOR2X1 U320 ( .A(n387), .B(n389), .Y(n452) );
  XNOR2X1 U321 ( .A(n455), .B(n456), .Y(n176) );
  XOR2X1 U322 ( .A(n418), .B(n417), .Y(n419) );
  NAND2X1 U323 ( .A(n104), .B(b[9]), .Y(n444) );
  XNOR3X2 U324 ( .A(n409), .B(n362), .C(n361), .Y(n374) );
  XNOR2X1 U325 ( .A(n408), .B(n411), .Y(n361) );
  OAI2BB1X1 U326 ( .A0N(n87), .A1N(n167), .B0(n166), .Y(n168) );
  OAI21XL U327 ( .A0(n165), .A1(n182), .B0(n92), .Y(n166) );
  INVX1 U328 ( .A(n92), .Y(n164) );
  NAND2BX1 U329 ( .AN(n61), .B(n39), .Y(n383) );
  XNOR3X2 U330 ( .A(n80), .B(n81), .C(n396), .Y(n131) );
  XOR3X2 U331 ( .A(n136), .B(n135), .C(n134), .Y(n137) );
  XOR2X1 U332 ( .A(n443), .B(n442), .Y(n447) );
  NOR2X1 U333 ( .A(n387), .B(n490), .Y(n442) );
  AOI22X1 U334 ( .A0(n25), .A1(n441), .B0(n23), .B1(n440), .Y(n443) );
  OAI21XL U335 ( .A0(n23), .A1(n378), .B0(n60), .Y(n441) );
  OAI2BB1X1 U336 ( .A0N(n28), .A1N(n251), .B0(n250), .Y(n252) );
  AOI21X1 U337 ( .A0(n96), .A1(n217), .B0(n216), .Y(n219) );
  XOR3X2 U338 ( .A(n179), .B(n178), .C(n177), .Y(n189) );
  XOR2X1 U339 ( .A(n384), .B(n416), .Y(n420) );
  XOR2X1 U340 ( .A(n394), .B(n415), .Y(n422) );
  XOR2X1 U341 ( .A(n414), .B(n413), .Y(n415) );
  XOR3X2 U342 ( .A(n412), .B(n376), .C(n375), .Y(n394) );
  XOR2X1 U343 ( .A(n480), .B(n479), .Y(n481) );
  XOR2X1 U344 ( .A(n478), .B(n477), .Y(n479) );
  XOR2X1 U345 ( .A(n476), .B(n475), .Y(n480) );
  NOR2BX1 U346 ( .AN(n39), .B(n34), .Y(n298) );
  NOR2BX1 U347 ( .AN(a[12]), .B(n87), .Y(n143) );
  OAI21XL U348 ( .A0(n187), .A1(n182), .B0(n95), .Y(n188) );
  NOR2BX1 U349 ( .AN(n39), .B(n28), .Y(n249) );
  NOR2BX1 U350 ( .AN(n39), .B(n86), .Y(n128) );
  XNOR3X2 U351 ( .A(n347), .B(n346), .C(n343), .Y(n348) );
  XOR3X2 U352 ( .A(n339), .B(n338), .C(n337), .Y(n343) );
  XOR2X1 U353 ( .A(n385), .B(n501), .Y(n347) );
  NAND2BXL U354 ( .AN(n97), .B(n39), .Y(n226) );
  AND2X2 U355 ( .A(n11), .B(a[3]), .Y(n155) );
  XNOR3X2 U356 ( .A(n82), .B(n83), .C(n436), .Y(n146) );
  AND2X2 U357 ( .A(n37), .B(n95), .Y(n170) );
  NAND2BXL U358 ( .AN(b[9]), .B(n47), .Y(n317) );
  XNOR2X1 U359 ( .A(n438), .B(n435), .Y(n151) );
  XNOR2X1 U360 ( .A(n450), .B(n451), .Y(n193) );
  XNOR2X1 U361 ( .A(n330), .B(n329), .Y(n331) );
  XOR2X1 U362 ( .A(n494), .B(n491), .Y(n329) );
  XNOR3X2 U363 ( .A(n327), .B(n493), .C(n362), .Y(n330) );
  INVX1 U364 ( .A(n98), .Y(n320) );
  OAI21XL U365 ( .A0(n20), .A1(n496), .B0(n8), .Y(n483) );
  NOR2X1 U366 ( .A(n490), .B(n495), .Y(n459) );
  INVX1 U367 ( .A(n101), .Y(n495) );
  XOR2X1 U368 ( .A(n306), .B(n305), .Y(n333) );
  NOR2X1 U369 ( .A(n387), .B(n49), .Y(n399) );
  XNOR3X2 U370 ( .A(n365), .B(n364), .C(n363), .Y(n373) );
  NAND2X1 U371 ( .A(n34), .B(a[1]), .Y(n352) );
  NAND2X1 U372 ( .A(n100), .B(n32), .Y(n353) );
  XOR2X1 U373 ( .A(n355), .B(n354), .Y(n356) );
  XOR2X1 U374 ( .A(n428), .B(n427), .Y(n429) );
  XOR2X1 U375 ( .A(n470), .B(n469), .Y(n471) );
  INVX1 U376 ( .A(n100), .Y(n387) );
  XOR2X1 U377 ( .A(n426), .B(n425), .Y(n430) );
  AOI22X1 U378 ( .A0(a[0]), .A1(n434), .B0(n25), .B1(n433), .Y(n439) );
  OAI21XL U379 ( .A0(n25), .A1(n496), .B0(n8), .Y(n434) );
  OAI21XL U380 ( .A0(n100), .A1(n49), .B0(n35), .Y(n433) );
  XOR2X1 U381 ( .A(n367), .B(n366), .Y(n368) );
  INVX1 U382 ( .A(b[0]), .Y(n497) );
  OAI2BB1X1 U383 ( .A0N(n86), .A1N(n130), .B0(n129), .Y(n132) );
  BUFX3 U384 ( .A(a[4]), .Y(n102) );
  BUFX3 U385 ( .A(a[6]), .Y(n104) );
  BUFX3 U386 ( .A(a[2]), .Y(n101) );
  BUFX3 U387 ( .A(a[5]), .Y(n103) );
  BUFX3 U388 ( .A(b[10]), .Y(n98) );
  BUFX3 U389 ( .A(b[11]), .Y(n99) );
  BUFX3 U390 ( .A(b[3]), .Y(n87) );
  BUFX3 U391 ( .A(b[4]), .Y(n92) );
  BUFX3 U392 ( .A(b[5]), .Y(n95) );
  BUFX3 U393 ( .A(b[6]), .Y(n96) );
  BUFX3 U394 ( .A(b[7]), .Y(n97) );
  INVX1 U395 ( .A(b[1]), .Y(n496) );
  BUFX3 U396 ( .A(a[0]), .Y(n100) );
  BUFX3 U397 ( .A(b[2]), .Y(n86) );
  OAI21XL U398 ( .A0(n111), .A1(n381), .B0(n26), .Y(n122) );
  OAI21XL U399 ( .A0(n180), .A1(n381), .B0(n92), .Y(n181) );
  OAI21XL U400 ( .A0(n298), .A1(n381), .B0(n28), .Y(n299) );
  AOI21XL U401 ( .A0(n316), .A1(n215), .B0(n214), .Y(n216) );
  OAI21XL U402 ( .A0(n128), .A1(n381), .B0(b[1]), .Y(n129) );
  AOI21XL U403 ( .A0(n316), .A1(n226), .B0(n225), .Y(n230) );
  OAI21XL U404 ( .A0(n249), .A1(n381), .B0(n97), .Y(n250) );
  AOI2BB2X1 U405 ( .B0(b[0]), .B1(n381), .A0N(n85), .A1N(n378), .Y(n382) );
  OAI2BB1XL U406 ( .A0N(a[12]), .A1N(n164), .B0(n316), .Y(n167) );
  NAND2BX4 U407 ( .AN(a[11]), .B(a[12]), .Y(n316) );
endmodule


module multiplier_10 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n36, n37, n38, n39, n43, n47, n49, n50, n51, n52,
         n53, n54, n55, n57, n58, n59, n61, n63, n64, n74, n77, n81, n83, n84,
         n85, n86, n87, n92, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n122, n127, n128,
         n131, n132, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n202, n203, n204, n205, n210,
         n211, n212, n213, n214, n215, n216, n217, n219, n220, n221, n239,
         n240, n246, n247, n248, n249, n250, n251, n252, n253, n254, n259,
         n260, n261, n262, n263, n264, n265, n266, n286, n288, n289, n290,
         n291, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n311, n314, n315, n316, n317, n318, n319, n320, n321, n323,
         n324, n325, n326, n327, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531;

  NOR2XL U1 ( .A(n32), .B(n103), .Y(n169) );
  NOR2X1 U2 ( .A(n24), .B(n32), .Y(n298) );
  OAI221XL U3 ( .A0(n108), .A1(n58), .B0(n7), .B1(n32), .C0(n366), .Y(n367) );
  OAI2BB1X1 U4 ( .A0N(n26), .A1N(n34), .B0(n365), .Y(n300) );
  AND2X2 U5 ( .A(n84), .B(n102), .Y(n513) );
  NOR2X1 U6 ( .A(n32), .B(n85), .Y(n143) );
  OAI21XL U7 ( .A0(n1), .A1(n84), .B0(n365), .Y(n145) );
  INVXL U8 ( .A(n103), .Y(n1) );
  OAI21XL U9 ( .A0(n2), .A1(n92), .B0(n365), .Y(n219) );
  INVX1 U10 ( .A(n34), .Y(n2) );
  OAI21XL U11 ( .A0(b[10]), .A1(n32), .B0(n305), .Y(n315) );
  NOR2X1 U12 ( .A(n512), .B(n14), .Y(n404) );
  XNOR3X2 U13 ( .A(n374), .B(n458), .C(n180), .Y(c[2]) );
  BUFX4 U14 ( .A(b[3]), .Y(n85) );
  OAI21X1 U15 ( .A0(n372), .A1(n371), .B0(n370), .Y(n441) );
  INVX2 U16 ( .A(n142), .Y(n326) );
  XOR2X1 U17 ( .A(n457), .B(n456), .Y(n486) );
  XOR2X1 U18 ( .A(n107), .B(n63), .Y(n142) );
  NAND2BX2 U19 ( .AN(a[12]), .B(n103), .Y(n365) );
  CLKBUFX2 U20 ( .A(b[11]), .Y(n30) );
  AOI21X2 U21 ( .A0(n30), .A1(n106), .B0(n105), .Y(n107) );
  NAND2BX2 U22 ( .AN(n103), .B(a[12]), .Y(n305) );
  BUFX8 U23 ( .A(a[11]), .Y(n103) );
  OAI2BB1X1 U24 ( .A0N(n103), .A1N(n187), .B0(n365), .Y(n190) );
  NOR2X1 U25 ( .A(n259), .B(n254), .Y(n264) );
  NAND2BX1 U26 ( .AN(a[12]), .B(n34), .Y(n166) );
  INVX1 U27 ( .A(n32), .Y(n33) );
  INVX1 U28 ( .A(a[12]), .Y(n32) );
  INVX1 U29 ( .A(b[10]), .Y(n306) );
  BUFX3 U30 ( .A(a[11]), .Y(n34) );
  XNOR3X2 U31 ( .A(n54), .B(n55), .C(n301), .Y(n3) );
  INVX1 U32 ( .A(b[0]), .Y(n4) );
  INVX1 U33 ( .A(n383), .Y(n5) );
  BUFX3 U34 ( .A(n58), .Y(n6) );
  NAND2X1 U35 ( .A(b[1]), .B(n525), .Y(n58) );
  NAND2X1 U36 ( .A(b[0]), .B(n524), .Y(n7) );
  NAND2X1 U37 ( .A(b[0]), .B(n524), .Y(n57) );
  INVX1 U38 ( .A(n187), .Y(n8) );
  INVX1 U39 ( .A(n86), .Y(n187) );
  INVX1 U40 ( .A(n306), .Y(n9) );
  INVX1 U41 ( .A(n384), .Y(n10) );
  INVX1 U42 ( .A(n382), .Y(n11) );
  INVX1 U43 ( .A(a[10]), .Y(n12) );
  INVX1 U44 ( .A(n12), .Y(n13) );
  INVX1 U45 ( .A(a[9]), .Y(n14) );
  INVX1 U46 ( .A(n14), .Y(n15) );
  INVX1 U47 ( .A(n14), .Y(n16) );
  INVX1 U48 ( .A(a[8]), .Y(n17) );
  INVX1 U49 ( .A(n17), .Y(n18) );
  INVX1 U50 ( .A(a[7]), .Y(n19) );
  INVXL U51 ( .A(n19), .Y(n20) );
  INVX1 U52 ( .A(n455), .Y(n21) );
  INVX1 U53 ( .A(n523), .Y(n22) );
  INVX1 U54 ( .A(b[9]), .Y(n23) );
  INVX1 U55 ( .A(n23), .Y(n24) );
  INVX1 U56 ( .A(n23), .Y(n25) );
  INVX1 U57 ( .A(b[8]), .Y(n26) );
  INVX1 U58 ( .A(n26), .Y(n27) );
  INVXL U59 ( .A(n26), .Y(n28) );
  INVX1 U60 ( .A(n251), .Y(n29) );
  INVX2 U61 ( .A(n486), .Y(n376) );
  OAI21XL U62 ( .A0(n102), .A1(n364), .B0(n58), .Y(n491) );
  XOR2X2 U63 ( .A(n141), .B(n140), .Y(n178) );
  XOR2X2 U64 ( .A(n39), .B(n177), .Y(n38) );
  NOR2X2 U65 ( .A(n368), .B(n384), .Y(n369) );
  BUFX3 U66 ( .A(b[4]), .Y(n31) );
  NAND2BXL U67 ( .AN(n92), .B(n33), .Y(n252) );
  OAI2BB1X2 U68 ( .A0N(n34), .A1N(n306), .B0(n365), .Y(n106) );
  OAI2BB1XL U69 ( .A0N(n103), .A1N(b[4]), .B0(n384), .Y(n370) );
  INVX1 U70 ( .A(n305), .Y(n371) );
  XOR2X1 U71 ( .A(n485), .B(n484), .Y(c[5]) );
  XNOR2X1 U72 ( .A(n326), .B(n64), .Y(n363) );
  NAND2BXL U73 ( .AN(b[11]), .B(a[12]), .Y(n104) );
  NAND2BXL U74 ( .AN(n87), .B(n33), .Y(n188) );
  XNOR2X1 U75 ( .A(n297), .B(n296), .Y(n55) );
  XNOR2X1 U76 ( .A(n291), .B(n36), .Y(n59) );
  AOI21X1 U77 ( .A0(n87), .A1(n190), .B0(n189), .Y(n205) );
  XNOR2X1 U78 ( .A(n373), .B(n36), .Y(n51) );
  AOI22X1 U79 ( .A0(n20), .A1(n511), .B0(n18), .B1(n510), .Y(n514) );
  NAND2XL U80 ( .A(a[8]), .B(n86), .Y(n81) );
  NAND2XL U81 ( .A(n85), .B(n102), .Y(n530) );
  NOR2BX1 U82 ( .AN(n103), .B(n25), .Y(n311) );
  INVXL U83 ( .A(n286), .Y(n214) );
  INVXL U84 ( .A(n363), .Y(n179) );
  XOR3X2 U85 ( .A(n37), .B(n264), .C(n263), .Y(n36) );
  XNOR2X1 U86 ( .A(n250), .B(n249), .Y(n37) );
  XOR3X2 U87 ( .A(n459), .B(n460), .C(n163), .Y(n39) );
  NOR2XL U88 ( .A(n378), .B(n383), .Y(n408) );
  INVXL U89 ( .A(n377), .Y(n373) );
  XOR2XL U90 ( .A(n291), .B(n3), .Y(n332) );
  NOR2XL U91 ( .A(n381), .B(n384), .Y(n463) );
  NOR2XL U92 ( .A(n380), .B(n383), .Y(n506) );
  XNOR2X1 U93 ( .A(n486), .B(n375), .Y(n180) );
  XOR3X2 U94 ( .A(n43), .B(n395), .C(n47), .Y(n347) );
  XOR3X2 U95 ( .A(n396), .B(n334), .C(n333), .Y(n43) );
  XNOR3X2 U96 ( .A(n346), .B(n339), .C(n338), .Y(n47) );
  XOR2X1 U97 ( .A(n61), .B(n436), .Y(c[1]) );
  INVXL U98 ( .A(n103), .Y(n108) );
  AOI22XL U99 ( .A0(n11), .A1(n110), .B0(n30), .B1(n109), .Y(n375) );
  NAND2XL U100 ( .A(n92), .B(n102), .Y(n387) );
  INVXL U101 ( .A(n84), .Y(n512) );
  AOI21XL U102 ( .A0(n34), .A1(n167), .B0(n368), .Y(n173) );
  INVXL U103 ( .A(b[4]), .Y(n167) );
  AOI22XL U104 ( .A0(n98), .A1(n465), .B0(n99), .B1(n464), .Y(n467) );
  NAND2XL U105 ( .A(n25), .B(a[10]), .Y(n221) );
  NAND2XL U106 ( .A(n5), .B(n99), .Y(n334) );
  NAND2XL U107 ( .A(a[7]), .B(n25), .Y(n460) );
  NAND2XL U108 ( .A(n92), .B(n18), .Y(n443) );
  AOI22XL U109 ( .A0(n18), .A1(n527), .B0(n16), .B1(n526), .Y(n528) );
  NAND2XL U110 ( .A(n27), .B(a[8]), .Y(n165) );
  NAND2XL U111 ( .A(n92), .B(n15), .Y(n164) );
  NAND2XL U112 ( .A(n100), .B(n24), .Y(n389) );
  NAND2XL U113 ( .A(n101), .B(n27), .Y(n391) );
  NAND2XL U114 ( .A(n95), .B(n98), .Y(n150) );
  NAND2XL U115 ( .A(n99), .B(b[11]), .Y(n149) );
  INVXL U116 ( .A(n92), .Y(n383) );
  NAND2XL U117 ( .A(a[10]), .B(n95), .Y(n63) );
  NAND2XL U118 ( .A(n20), .B(n11), .Y(n246) );
  NAND2XL U119 ( .A(n18), .B(n9), .Y(n260) );
  XNOR3X2 U120 ( .A(n49), .B(n401), .C(n316), .Y(n531) );
  NAND2XL U121 ( .A(n16), .B(n95), .Y(n49) );
  OAI2BB1X1 U122 ( .A0N(n85), .A1N(n145), .B0(n144), .Y(n147) );
  NAND2XL U123 ( .A(n31), .B(n20), .Y(n406) );
  NAND2XL U124 ( .A(n31), .B(n101), .Y(n529) );
  NAND2XL U125 ( .A(n96), .B(n25), .Y(n324) );
  NAND2XL U126 ( .A(n92), .B(n98), .Y(n323) );
  NAND2XL U127 ( .A(n84), .B(n13), .Y(n412) );
  NAND2XL U128 ( .A(n13), .B(n85), .Y(n139) );
  NAND2XL U129 ( .A(n99), .B(n31), .Y(n504) );
  NAND2XL U130 ( .A(n102), .B(n9), .Y(n459) );
  INVXL U131 ( .A(n101), .Y(n378) );
  NAND2XL U132 ( .A(n87), .B(a[6]), .Y(n409) );
  NAND2XL U133 ( .A(n21), .B(n86), .Y(n508) );
  NAND2XL U134 ( .A(n29), .B(n98), .Y(n507) );
  NAND2XL U135 ( .A(n31), .B(n18), .Y(n413) );
  NAND2XL U136 ( .A(n102), .B(n24), .Y(n447) );
  NAND2XL U137 ( .A(n21), .B(n28), .Y(n400) );
  NAND2XL U138 ( .A(n28), .B(n97), .Y(n317) );
  NAND2XL U139 ( .A(n96), .B(n5), .Y(n289) );
  NAND2XL U140 ( .A(n102), .B(b[11]), .Y(n473) );
  NAND2XL U141 ( .A(n29), .B(n96), .Y(n487) );
  NAND2XL U142 ( .A(n100), .B(n31), .Y(n515) );
  NAND2XL U143 ( .A(n100), .B(b[11]), .Y(n449) );
  NAND2XL U144 ( .A(n15), .B(n30), .Y(n296) );
  NAND2XL U145 ( .A(n18), .B(b[11]), .Y(n240) );
  NOR2BXL U146 ( .AN(n33), .B(n28), .Y(n216) );
  XOR2X1 U147 ( .A(n202), .B(n195), .Y(n203) );
  NOR2BXL U148 ( .AN(a[12]), .B(n86), .Y(n168) );
  NAND2XL U149 ( .A(n86), .B(n13), .Y(n442) );
  NAND2XL U150 ( .A(a[8]), .B(n95), .Y(n297) );
  NAND2XL U151 ( .A(n101), .B(n95), .Y(n194) );
  NAND2XL U152 ( .A(n24), .B(a[8]), .Y(n193) );
  NAND2XL U153 ( .A(n100), .B(n95), .Y(n461) );
  NAND2XL U154 ( .A(n101), .B(n30), .Y(n462) );
  NAND2XL U155 ( .A(n87), .B(n99), .Y(n318) );
  INVXL U156 ( .A(n99), .Y(n455) );
  NAND2XL U157 ( .A(n22), .B(n25), .Y(n399) );
  NAND2XL U158 ( .A(n86), .B(n97), .Y(n488) );
  NAND2XL U159 ( .A(n101), .B(n85), .Y(n516) );
  NAND2XL U160 ( .A(a[7]), .B(n9), .Y(n474) );
  NAND2XL U161 ( .A(n101), .B(n9), .Y(n450) );
  NAND2XL U162 ( .A(n100), .B(n29), .Y(n335) );
  NAND2XL U163 ( .A(n25), .B(n97), .Y(n337) );
  NAND2XL U164 ( .A(n87), .B(a[7]), .Y(n388) );
  NAND2XL U165 ( .A(n92), .B(n20), .Y(n433) );
  NAND2XL U166 ( .A(n85), .B(n20), .Y(n398) );
  NAND2XL U167 ( .A(n31), .B(a[6]), .Y(n397) );
  NAND2XL U168 ( .A(a[5]), .B(n86), .Y(n333) );
  NAND2XL U169 ( .A(n85), .B(n16), .Y(n414) );
  NAND2XL U170 ( .A(a[7]), .B(n28), .Y(n448) );
  NAND2XL U171 ( .A(n99), .B(n85), .Y(n496) );
  NAND2XL U172 ( .A(n98), .B(n31), .Y(n495) );
  NAND2XL U173 ( .A(n92), .B(a[10]), .Y(n192) );
  NAND2XL U174 ( .A(n27), .B(n16), .Y(n191) );
  AOI22XL U175 ( .A0(n13), .A1(n403), .B0(n34), .B1(n402), .Y(n405) );
  NAND2XL U176 ( .A(n10), .B(n18), .Y(n407) );
  XNOR2X1 U177 ( .A(n50), .B(n319), .Y(n320) );
  NAND2XL U178 ( .A(n20), .B(n84), .Y(n50) );
  XOR3X2 U179 ( .A(n376), .B(n51), .C(n52), .Y(n484) );
  XNOR3X2 U180 ( .A(n375), .B(n483), .C(n374), .Y(n52) );
  XOR3X2 U181 ( .A(n53), .B(n302), .C(n332), .Y(n303) );
  NAND2XL U182 ( .A(n29), .B(n97), .Y(n53) );
  AOI22XL U183 ( .A0(a[6]), .A1(n501), .B0(n20), .B1(n500), .Y(n503) );
  NAND2XL U184 ( .A(n100), .B(n85), .Y(n505) );
  XNOR3X2 U185 ( .A(n327), .B(n326), .C(n528), .Y(n330) );
  NAND2XL U186 ( .A(n96), .B(n31), .Y(n212) );
  AOI22XL U187 ( .A0(n21), .A1(n470), .B0(a[4]), .B1(n469), .Y(n472) );
  NAND2XL U188 ( .A(n95), .B(n97), .Y(n111) );
  NAND2XL U189 ( .A(b[11]), .B(n98), .Y(n122) );
  NAND2XL U190 ( .A(n87), .B(a[8]), .Y(n74) );
  NAND2XL U191 ( .A(n15), .B(n86), .Y(n77) );
  NAND2XL U192 ( .A(n15), .B(b[4]), .Y(n83) );
  INVXL U193 ( .A(n100), .Y(n492) );
  NAND2XL U194 ( .A(n96), .B(n11), .Y(n419) );
  NAND2XL U195 ( .A(n86), .B(n20), .Y(n410) );
  NAND2XL U196 ( .A(n30), .B(n13), .Y(n401) );
  AND2X1 U197 ( .A(n33), .B(n95), .Y(n64) );
  NAND2XL U198 ( .A(n101), .B(n25), .Y(n435) );
  NAND2XL U199 ( .A(n102), .B(n28), .Y(n432) );
  INVXL U200 ( .A(n95), .Y(n382) );
  AND2X1 U201 ( .A(n13), .B(b[4]), .Y(n148) );
  AND2X1 U202 ( .A(n87), .B(a[10]), .Y(n176) );
  AND2X1 U203 ( .A(n16), .B(b[10]), .Y(n239) );
  AND2X1 U204 ( .A(n100), .B(n86), .Y(n319) );
  NAND2XL U205 ( .A(n13), .B(n9), .Y(n54) );
  XOR2X1 U206 ( .A(n446), .B(n445), .Y(n454) );
  XOR2X1 U207 ( .A(n444), .B(n443), .Y(n445) );
  NAND2XL U208 ( .A(n87), .B(n16), .Y(n444) );
  INVX2 U209 ( .A(n85), .Y(n384) );
  INVX1 U210 ( .A(n166), .Y(n368) );
  NAND2XL U211 ( .A(n28), .B(n98), .Y(n339) );
  NAND2XL U212 ( .A(n96), .B(n30), .Y(n356) );
  NAND2XL U213 ( .A(a[6]), .B(n8), .Y(n352) );
  NAND2XL U214 ( .A(a[5]), .B(n29), .Y(n353) );
  NAND2XL U215 ( .A(a[4]), .B(n5), .Y(n354) );
  NAND2XL U216 ( .A(n21), .B(n25), .Y(n422) );
  NAND2XL U217 ( .A(n31), .B(a[1]), .Y(n479) );
  NAND2XL U218 ( .A(n97), .B(n30), .Y(n424) );
  AND2X1 U219 ( .A(n18), .B(n84), .Y(n395) );
  AND2X1 U220 ( .A(n28), .B(a[0]), .Y(n521) );
  NAND2XL U221 ( .A(n10), .B(n97), .Y(n210) );
  NAND2XL U222 ( .A(n21), .B(n84), .Y(n478) );
  NAND2XL U223 ( .A(a[4]), .B(n28), .Y(n423) );
  AOI2BB2XL U224 ( .B0(b[0]), .B1(n371), .A0N(n365), .A1N(n364), .Y(n366) );
  INVXL U225 ( .A(b[1]), .Y(n364) );
  NAND2BXL U226 ( .AN(b[1]), .B(n34), .Y(n132) );
  XNOR2X1 U227 ( .A(n38), .B(n373), .Y(n286) );
  XOR2X1 U228 ( .A(n59), .B(n376), .Y(n265) );
  INVX1 U229 ( .A(n332), .Y(n348) );
  XNOR3X2 U230 ( .A(n349), .B(n348), .C(n347), .Y(c[10]) );
  XOR2X1 U231 ( .A(n142), .B(n375), .Y(n349) );
  XOR2X1 U232 ( .A(n531), .B(n3), .Y(n351) );
  XOR3X2 U233 ( .A(n262), .B(n261), .C(n260), .Y(n263) );
  XOR3X2 U234 ( .A(n351), .B(n521), .C(n522), .Y(c[8]) );
  XNOR3X2 U235 ( .A(n179), .B(n38), .C(n178), .Y(n181) );
  XOR3X2 U236 ( .A(n506), .B(n36), .C(n377), .Y(n385) );
  XNOR3X2 U237 ( .A(n38), .B(n499), .C(n215), .Y(n266) );
  XOR2X1 U238 ( .A(n489), .B(n64), .Y(n215) );
  XOR2X1 U239 ( .A(n498), .B(n497), .Y(n499) );
  XOR2X1 U240 ( .A(n488), .B(n487), .Y(n489) );
  XOR3X2 U241 ( .A(n359), .B(n358), .C(n357), .Y(n360) );
  XOR2X1 U242 ( .A(n399), .B(n400), .Y(n358) );
  XNOR3X2 U243 ( .A(n406), .B(n356), .C(n355), .Y(n357) );
  XOR2X1 U244 ( .A(n375), .B(n64), .Y(n359) );
  XNOR3X2 U245 ( .A(n176), .B(n175), .C(n174), .Y(n177) );
  XOR2X1 U246 ( .A(n266), .B(n265), .Y(c[6]) );
  XOR2X1 U247 ( .A(n429), .B(n428), .Y(c[12]) );
  XOR2X1 U248 ( .A(n520), .B(n519), .Y(n522) );
  XOR2X1 U249 ( .A(n518), .B(n517), .Y(n519) );
  XOR2X1 U250 ( .A(n385), .B(n509), .Y(n520) );
  XOR2X1 U251 ( .A(n516), .B(n515), .Y(n517) );
  XOR2X1 U252 ( .A(n468), .B(n463), .Y(n182) );
  XOR2X1 U253 ( .A(n467), .B(n466), .Y(n468) );
  NOR2X1 U254 ( .A(n380), .B(n512), .Y(n466) );
  XOR3X2 U255 ( .A(n179), .B(n178), .C(n374), .Y(n61) );
  XNOR3X2 U256 ( .A(n61), .B(n214), .C(n213), .Y(c[4]) );
  XNOR2X1 U257 ( .A(n304), .B(n303), .Y(c[7]) );
  XOR3X2 U258 ( .A(n182), .B(n181), .C(n180), .Y(c[3]) );
  XNOR3X2 U259 ( .A(n331), .B(n59), .C(n330), .Y(c[9]) );
  XNOR3X2 U260 ( .A(n362), .B(n361), .C(n360), .Y(c[11]) );
  NOR2X1 U261 ( .A(n512), .B(n378), .Y(n502) );
  OAI21XL U262 ( .A0(n30), .A1(n108), .B0(n365), .Y(n110) );
  OAI21XL U263 ( .A0(n16), .A1(n524), .B0(n6), .Y(n527) );
  OAI21XL U264 ( .A0(n18), .A1(n4), .B0(n57), .Y(n526) );
  OAI21XL U265 ( .A0(n311), .A1(n368), .B0(n9), .Y(n314) );
  OAI21XL U266 ( .A0(n99), .A1(n364), .B0(n58), .Y(n465) );
  OAI21XL U267 ( .A0(n98), .A1(n4), .B0(n57), .Y(n464) );
  AOI22X1 U268 ( .A0(n13), .A1(n394), .B0(n16), .B1(n393), .Y(n396) );
  OAI21XL U269 ( .A0(n13), .A1(n364), .B0(n58), .Y(n393) );
  OAI21XL U270 ( .A0(n16), .A1(n4), .B0(n57), .Y(n394) );
  INVXL U271 ( .A(n87), .Y(n251) );
  OAI2BB1X1 U272 ( .A0N(n25), .A1N(n315), .B0(n314), .Y(n316) );
  OAI21XL U273 ( .A0(n18), .A1(n364), .B0(n58), .Y(n511) );
  OAI21XL U274 ( .A0(n100), .A1(n364), .B0(n58), .Y(n470) );
  OAI21XL U275 ( .A0(n20), .A1(n364), .B0(n58), .Y(n501) );
  OAI21XL U276 ( .A0(n103), .A1(n364), .B0(n58), .Y(n403) );
  OAI21XL U277 ( .A0(n101), .A1(n4), .B0(n57), .Y(n490) );
  OAI21XL U278 ( .A0(n20), .A1(n4), .B0(n7), .Y(n510) );
  OAI21XL U279 ( .A0(n97), .A1(n525), .B0(n57), .Y(n437) );
  OAI21XL U280 ( .A0(n99), .A1(n4), .B0(n7), .Y(n469) );
  AOI22X1 U281 ( .A0(a[4]), .A1(n476), .B0(a[5]), .B1(n475), .Y(n477) );
  OAI21XL U282 ( .A0(a[5]), .A1(n364), .B0(n6), .Y(n476) );
  OAI21XL U283 ( .A0(a[4]), .A1(n525), .B0(n7), .Y(n475) );
  OAI21XL U284 ( .A0(a[6]), .A1(n4), .B0(n57), .Y(n500) );
  OAI21XL U285 ( .A0(n13), .A1(n4), .B0(n7), .Y(n402) );
  OAI21XL U286 ( .A0(n173), .A1(n187), .B0(n170), .Y(n174) );
  OAI21XL U287 ( .A0(n169), .A1(n168), .B0(n31), .Y(n170) );
  MXI2X1 U288 ( .A(n32), .B(n369), .S0(b[4]), .Y(n372) );
  XOR2X1 U289 ( .A(n162), .B(n153), .Y(n374) );
  XNOR3X2 U290 ( .A(n434), .B(n152), .C(n151), .Y(n153) );
  XNOR3X2 U291 ( .A(n148), .B(n147), .C(n146), .Y(n162) );
  NAND2X1 U292 ( .A(n100), .B(n9), .Y(n434) );
  XNOR3X2 U293 ( .A(n387), .B(n131), .C(n128), .Y(n141) );
  XNOR3X2 U294 ( .A(n139), .B(n138), .C(n137), .Y(n140) );
  XNOR3X2 U295 ( .A(n205), .B(n204), .C(n203), .Y(n377) );
  XNOR2X1 U296 ( .A(n474), .B(n473), .Y(n204) );
  XOR2X1 U297 ( .A(n248), .B(n247), .Y(n291) );
  XOR2X1 U298 ( .A(n246), .B(n240), .Y(n247) );
  XNOR3X2 U299 ( .A(n239), .B(n221), .C(n220), .Y(n248) );
  NOR2X1 U300 ( .A(n382), .B(n455), .Y(n456) );
  XOR2X1 U301 ( .A(n454), .B(n453), .Y(n457) );
  NAND2X1 U302 ( .A(n102), .B(n95), .Y(n261) );
  NOR2BX1 U303 ( .AN(a[12]), .B(n84), .Y(n134) );
  NAND2X1 U304 ( .A(a[7]), .B(n30), .Y(n249) );
  XOR2X1 U305 ( .A(n150), .B(n149), .Y(n152) );
  OAI21XL U306 ( .A0(n143), .A1(n371), .B0(n84), .Y(n144) );
  XOR2X1 U307 ( .A(n496), .B(n495), .Y(n497) );
  XNOR2X1 U308 ( .A(n192), .B(n191), .Y(n202) );
  AND2X2 U309 ( .A(n8), .B(n96), .Y(n483) );
  XNOR3X2 U310 ( .A(n392), .B(n349), .C(n178), .Y(c[0]) );
  NOR2X1 U311 ( .A(n381), .B(n4), .Y(n392) );
  XOR2X1 U312 ( .A(n290), .B(n289), .Y(n302) );
  NAND2X1 U313 ( .A(n8), .B(n98), .Y(n290) );
  XOR2X1 U314 ( .A(n440), .B(n439), .Y(n458) );
  NOR2X1 U315 ( .A(n381), .B(n512), .Y(n439) );
  AOI22X1 U316 ( .A0(n97), .A1(n438), .B0(n22), .B1(n437), .Y(n440) );
  OAI21XL U317 ( .A0(n22), .A1(n364), .B0(n58), .Y(n438) );
  XOR2X1 U318 ( .A(n165), .B(n164), .Y(n175) );
  XOR2X1 U319 ( .A(n389), .B(n391), .Y(n131) );
  XOR2X1 U320 ( .A(n194), .B(n193), .Y(n195) );
  XOR2X1 U321 ( .A(n452), .B(n451), .Y(n453) );
  XOR2X1 U322 ( .A(n448), .B(n447), .Y(n452) );
  XOR2X1 U323 ( .A(n450), .B(n449), .Y(n451) );
  XOR2X1 U324 ( .A(n416), .B(n415), .Y(n417) );
  XOR2X1 U325 ( .A(n414), .B(n413), .Y(n415) );
  XOR2X1 U326 ( .A(n367), .B(n412), .Y(n416) );
  XNOR3X2 U327 ( .A(n503), .B(n288), .C(n286), .Y(n304) );
  XOR3X2 U328 ( .A(n504), .B(n505), .C(n502), .Y(n288) );
  XNOR3X2 U329 ( .A(n405), .B(n351), .C(n350), .Y(n362) );
  XNOR2X1 U330 ( .A(n404), .B(n407), .Y(n350) );
  NAND2X1 U331 ( .A(n27), .B(a[10]), .Y(n250) );
  XNOR3X2 U332 ( .A(n321), .B(n320), .C(n531), .Y(n331) );
  XOR2X1 U333 ( .A(n318), .B(n317), .Y(n321) );
  OAI2BB1X1 U334 ( .A0N(n25), .A1N(n300), .B0(n299), .Y(n301) );
  OAI21XL U335 ( .A0(n298), .A1(n371), .B0(n28), .Y(n299) );
  XNOR3X2 U336 ( .A(n74), .B(n77), .C(n433), .Y(n146) );
  XNOR3X2 U337 ( .A(n81), .B(n83), .C(n388), .Y(n137) );
  XOR3X2 U338 ( .A(n529), .B(n530), .C(n325), .Y(n327) );
  XNOR3X2 U339 ( .A(n472), .B(n212), .C(n211), .Y(n213) );
  XOR2X1 U340 ( .A(n210), .B(n471), .Y(n211) );
  XNOR3X2 U341 ( .A(n127), .B(n122), .C(n111), .Y(n128) );
  NAND2X1 U342 ( .A(b[10]), .B(n99), .Y(n127) );
  NAND2X1 U343 ( .A(n24), .B(n15), .Y(n262) );
  OAI2BB1X1 U344 ( .A0N(n28), .A1N(n219), .B0(n217), .Y(n220) );
  OAI21XL U345 ( .A0(n216), .A1(n371), .B0(n92), .Y(n217) );
  XOR2X1 U346 ( .A(n494), .B(n493), .Y(n498) );
  NOR2X1 U347 ( .A(n512), .B(n492), .Y(n493) );
  AOI22X1 U348 ( .A0(n101), .A1(n491), .B0(n102), .B1(n490), .Y(n494) );
  XOR2X1 U349 ( .A(n514), .B(n513), .Y(n518) );
  XOR2X1 U350 ( .A(n421), .B(n420), .Y(n429) );
  XNOR2X1 U351 ( .A(n419), .B(n531), .Y(n420) );
  XOR2X1 U352 ( .A(n418), .B(n417), .Y(n421) );
  XOR2X1 U353 ( .A(n442), .B(n441), .Y(n446) );
  XOR2X1 U354 ( .A(n386), .B(n411), .Y(n418) );
  XOR2X1 U355 ( .A(n410), .B(n409), .Y(n411) );
  XOR2X1 U356 ( .A(n363), .B(n408), .Y(n386) );
  XOR2X1 U357 ( .A(n482), .B(n481), .Y(n485) );
  XOR2X1 U358 ( .A(n480), .B(n479), .Y(n481) );
  XOR2X1 U359 ( .A(n478), .B(n477), .Y(n482) );
  NAND2X1 U360 ( .A(n22), .B(n10), .Y(n480) );
  NAND2BX1 U361 ( .AN(n87), .B(n34), .Y(n253) );
  XNOR2X1 U362 ( .A(n435), .B(n432), .Y(n151) );
  XOR2X1 U363 ( .A(n461), .B(n462), .Y(n163) );
  AOI22X1 U364 ( .A0(a[0]), .A1(n431), .B0(a[1]), .B1(n430), .Y(n436) );
  OAI21XL U365 ( .A0(a[1]), .A1(n524), .B0(n6), .Y(n431) );
  OAI21XL U366 ( .A0(n96), .A1(n4), .B0(n7), .Y(n430) );
  NOR2X1 U367 ( .A(n512), .B(n523), .Y(n471) );
  INVX1 U368 ( .A(n98), .Y(n523) );
  XOR2X1 U369 ( .A(n508), .B(n507), .Y(n509) );
  XOR2X1 U370 ( .A(n427), .B(n426), .Y(n428) );
  XOR2X1 U371 ( .A(n423), .B(n422), .Y(n427) );
  XOR2X1 U372 ( .A(n425), .B(n424), .Y(n426) );
  NAND2X1 U373 ( .A(n22), .B(n9), .Y(n425) );
  XOR3X2 U374 ( .A(n337), .B(n336), .C(n335), .Y(n338) );
  NAND2X1 U375 ( .A(n96), .B(n9), .Y(n336) );
  XNOR3X2 U376 ( .A(n354), .B(n353), .C(n352), .Y(n361) );
  INVX1 U377 ( .A(n96), .Y(n381) );
  NAND2X1 U378 ( .A(a[1]), .B(n9), .Y(n355) );
  XOR2X1 U379 ( .A(n324), .B(n323), .Y(n325) );
  XOR2X1 U380 ( .A(n398), .B(n397), .Y(n346) );
  INVX1 U381 ( .A(n97), .Y(n380) );
  OAI2BB1X1 U382 ( .A0N(n84), .A1N(n136), .B0(n135), .Y(n138) );
  OAI21XL U383 ( .A0(n134), .A1(n371), .B0(b[1]), .Y(n135) );
  BUFX3 U384 ( .A(a[3]), .Y(n99) );
  BUFX3 U385 ( .A(a[6]), .Y(n102) );
  BUFX3 U386 ( .A(a[2]), .Y(n98) );
  BUFX3 U387 ( .A(a[4]), .Y(n100) );
  BUFX3 U388 ( .A(a[5]), .Y(n101) );
  BUFX3 U389 ( .A(a[1]), .Y(n97) );
  BUFX3 U390 ( .A(b[6]), .Y(n87) );
  BUFX3 U391 ( .A(b[12]), .Y(n95) );
  BUFX3 U392 ( .A(b[7]), .Y(n92) );
  INVX1 U393 ( .A(b[0]), .Y(n525) );
  INVX1 U394 ( .A(b[1]), .Y(n524) );
  BUFX3 U395 ( .A(b[5]), .Y(n86) );
  BUFX3 U396 ( .A(b[2]), .Y(n84) );
  BUFX3 U397 ( .A(a[0]), .Y(n96) );
  NAND2X1 U398 ( .A(n365), .B(n132), .Y(n136) );
  AOI21X1 U399 ( .A0(n365), .A1(n253), .B0(n383), .Y(n254) );
  OAI21XL U400 ( .A0(n11), .A1(n32), .B0(n305), .Y(n109) );
  AOI21X1 U401 ( .A0(n305), .A1(n188), .B0(n187), .Y(n189) );
  AOI21X1 U402 ( .A0(n305), .A1(n252), .B0(n251), .Y(n259) );
  AOI21X1 U403 ( .A0(n305), .A1(n104), .B0(n306), .Y(n105) );
endmodule


module multiplier_9 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n47, n49, n50, n51, n52,
         n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n92, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n119, n122, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n202,
         n203, n204, n205, n210, n211, n212, n213, n214, n215, n216, n217,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n230,
         n233, n234, n235, n236, n237, n238, n239, n240, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n259, n260, n261, n262, n263,
         n264, n265, n266, n278, n286, n288, n289, n290, n291, n292, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n343, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508;

  XOR2X2 U1 ( .A(n427), .B(n426), .Y(n429) );
  INVX1 U2 ( .A(n327), .Y(n387) );
  NAND2BXL U3 ( .AN(n103), .B(n111), .Y(n3) );
  OAI21XL U4 ( .A0(n1), .A1(n98), .B0(n327), .Y(n174) );
  INVXL U5 ( .A(n111), .Y(n1) );
  NOR2BX1 U6 ( .AN(n106), .B(n495), .Y(n479) );
  OAI211X1 U7 ( .A0(n2), .A1(n65), .B0(n389), .C0(n388), .Y(n394) );
  INVX1 U8 ( .A(n33), .Y(n2) );
  OAI2BB1X1 U9 ( .A0N(n327), .A1N(n3), .B0(n102), .Y(n122) );
  AOI211X1 U10 ( .A0(n328), .A1(n34), .B0(n333), .C0(n37), .Y(n4) );
  INVX1 U11 ( .A(n4), .Y(n337) );
  NOR2X1 U12 ( .A(n25), .B(n495), .Y(n460) );
  NOR2X1 U13 ( .A(n39), .B(n9), .Y(n127) );
  NAND3X1 U14 ( .A(n191), .B(n193), .C(n195), .Y(n204) );
  XOR3X2 U15 ( .A(n380), .B(n415), .C(n378), .Y(n381) );
  NAND3BX1 U16 ( .AN(n331), .B(n330), .C(n332), .Y(n336) );
  XOR3X2 U17 ( .A(n322), .B(n497), .C(n321), .Y(n346) );
  XNOR2X1 U18 ( .A(n230), .B(n444), .Y(c[1]) );
  BUFX3 U19 ( .A(n386), .Y(n96) );
  INVX1 U20 ( .A(n96), .Y(n189) );
  XOR2X2 U21 ( .A(n128), .B(n127), .Y(n384) );
  XNOR3X2 U22 ( .A(n251), .B(n250), .C(n249), .Y(n5) );
  XNOR3X2 U23 ( .A(n53), .B(n54), .C(n315), .Y(n6) );
  NAND2XL U24 ( .A(b[0]), .B(n501), .Y(n7) );
  INVX1 U25 ( .A(b[0]), .Y(n8) );
  INVX1 U26 ( .A(b[12]), .Y(n9) );
  INVX1 U27 ( .A(n9), .Y(n10) );
  INVX1 U28 ( .A(n9), .Y(n11) );
  INVX1 U29 ( .A(n398), .Y(n12) );
  INVX1 U30 ( .A(n223), .Y(n13) );
  BUFX3 U31 ( .A(n111), .Y(n14) );
  NAND2BX2 U32 ( .AN(n110), .B(n111), .Y(n327) );
  BUFX3 U33 ( .A(a[12]), .Y(n111) );
  INVX1 U34 ( .A(n413), .Y(n15) );
  INVX1 U35 ( .A(a[8]), .Y(n16) );
  INVX1 U36 ( .A(n16), .Y(n17) );
  INVX1 U37 ( .A(n16), .Y(n18) );
  INVX1 U38 ( .A(a[7]), .Y(n19) );
  INVXL U39 ( .A(n19), .Y(n20) );
  INVX1 U40 ( .A(n494), .Y(n21) );
  INVX1 U41 ( .A(a[3]), .Y(n22) );
  INVXL U42 ( .A(n22), .Y(n23) );
  INVX1 U43 ( .A(n500), .Y(n24) );
  INVX1 U44 ( .A(a[1]), .Y(n25) );
  INVX1 U45 ( .A(n25), .Y(n26) );
  INVX1 U46 ( .A(n129), .Y(n27) );
  OAI2BB1X2 U47 ( .A0N(n103), .A1N(n126), .B0(n122), .Y(n128) );
  INVX1 U48 ( .A(b[8]), .Y(n28) );
  INVX1 U49 ( .A(n28), .Y(n29) );
  INVXL U50 ( .A(n28), .Y(n30) );
  INVX1 U51 ( .A(n236), .Y(n31) );
  INVX1 U52 ( .A(n399), .Y(n32) );
  BUFX3 U53 ( .A(n110), .Y(n33) );
  INVX1 U54 ( .A(n119), .Y(n34) );
  INVX1 U55 ( .A(b[9]), .Y(n35) );
  INVX1 U56 ( .A(n35), .Y(n36) );
  INVXL U57 ( .A(n35), .Y(n37) );
  XOR2X2 U58 ( .A(n212), .B(n211), .Y(n290) );
  XNOR3X4 U59 ( .A(n178), .B(n51), .C(n52), .Y(n291) );
  XOR2X4 U60 ( .A(n291), .B(n179), .Y(n214) );
  NAND2BX2 U61 ( .AN(n111), .B(n110), .Y(n386) );
  INVX1 U62 ( .A(b[1]), .Y(n38) );
  INVX1 U63 ( .A(a[10]), .Y(n39) );
  INVX1 U64 ( .A(n39), .Y(n47) );
  INVXL U65 ( .A(n39), .Y(n49) );
  NAND2XL U66 ( .A(b[1]), .B(n502), .Y(n50) );
  XOR2X1 U67 ( .A(n290), .B(n79), .Y(n297) );
  BUFX3 U68 ( .A(a[11]), .Y(n110) );
  INVXL U69 ( .A(n333), .Y(n330) );
  NAND2BXL U70 ( .AN(n332), .B(n333), .Y(n334) );
  INVXL U71 ( .A(n384), .Y(n147) );
  NAND2X1 U72 ( .A(n100), .B(n109), .Y(n168) );
  NAND2X1 U73 ( .A(n101), .B(n17), .Y(n169) );
  NAND2X1 U74 ( .A(n47), .B(n103), .Y(n323) );
  XOR2XL U75 ( .A(n301), .B(n6), .Y(n369) );
  XNOR3X2 U76 ( .A(n167), .B(n451), .C(n84), .Y(n51) );
  XNOR3X2 U77 ( .A(n177), .B(n176), .C(n175), .Y(n52) );
  NAND2XL U78 ( .A(n196), .B(n194), .Y(n205) );
  XOR2X1 U79 ( .A(n82), .B(n452), .Y(c[2]) );
  NAND2XL U80 ( .A(n106), .B(n102), .Y(n442) );
  AOI22XL U81 ( .A0(n24), .A1(n459), .B0(n23), .B1(n458), .Y(n461) );
  AOI22XL U82 ( .A0(n18), .A1(n504), .B0(n15), .B1(n503), .Y(n506) );
  NAND2XL U83 ( .A(n101), .B(n108), .Y(n400) );
  AOI22XL U84 ( .A0(n49), .A1(n406), .B0(n15), .B1(n405), .Y(n407) );
  NAND2XL U85 ( .A(n96), .B(n148), .Y(n151) );
  NAND2XL U86 ( .A(n98), .B(n21), .Y(n408) );
  NAND2XL U87 ( .A(n107), .B(n102), .Y(n451) );
  NAND2XL U88 ( .A(n29), .B(n49), .Y(n247) );
  NAND2XL U89 ( .A(n36), .B(n49), .Y(n265) );
  NAND2BXL U90 ( .AN(n100), .B(n14), .Y(n224) );
  NAND2XL U91 ( .A(n109), .B(n10), .Y(n324) );
  NAND2XL U92 ( .A(n10), .B(n105), .Y(n162) );
  NAND2XL U93 ( .A(a[3]), .B(n103), .Y(n155) );
  NAND2XL U94 ( .A(n107), .B(n29), .Y(n403) );
  AOI22XL U95 ( .A0(n20), .A1(n493), .B0(n18), .B1(n492), .Y(n497) );
  AOI22XL U96 ( .A0(n49), .A1(n412), .B0(n33), .B1(n411), .Y(n415) );
  INVXL U97 ( .A(n100), .Y(n236) );
  NOR2X1 U98 ( .A(n240), .B(n239), .Y(n250) );
  AOI21XL U99 ( .A0(n96), .A1(n238), .B0(n398), .Y(n239) );
  NAND2XL U100 ( .A(n32), .B(n18), .Y(n417) );
  INVXL U101 ( .A(n109), .Y(n413) );
  NAND2XL U102 ( .A(n49), .B(n102), .Y(n53) );
  XNOR2X1 U103 ( .A(n303), .B(n302), .Y(n54) );
  NAND2XL U104 ( .A(n111), .B(n11), .Y(n373) );
  NAND2BXL U105 ( .AN(n102), .B(n14), .Y(n326) );
  NAND2XL U106 ( .A(n20), .B(n11), .Y(n286) );
  NAND2XL U107 ( .A(n96), .B(n304), .Y(n314) );
  NAND2XL U108 ( .A(n96), .B(n325), .Y(n328) );
  NAND2BXL U109 ( .AN(n36), .B(n33), .Y(n325) );
  NAND2XL U110 ( .A(n108), .B(n34), .Y(n453) );
  NAND2XL U111 ( .A(n36), .B(n109), .Y(n248) );
  NAND2XL U112 ( .A(n23), .B(b[4]), .Y(n490) );
  NAND2XL U113 ( .A(b[4]), .B(n26), .Y(n472) );
  INVXL U114 ( .A(n101), .Y(n398) );
  NAND2XL U115 ( .A(n107), .B(n11), .Y(n221) );
  NAND2XL U116 ( .A(n100), .B(n108), .Y(n419) );
  NAND2XL U117 ( .A(a[7]), .B(n102), .Y(n467) );
  NAND2XL U118 ( .A(n108), .B(n29), .Y(n440) );
  NAND2XL U119 ( .A(n107), .B(n36), .Y(n443) );
  NAND2XL U120 ( .A(n97), .B(n15), .Y(n423) );
  NAND2XL U121 ( .A(n98), .B(n18), .Y(n422) );
  NAND2XL U122 ( .A(n34), .B(n328), .Y(n332) );
  NAND2XL U123 ( .A(n109), .B(n103), .Y(n302) );
  NAND2XL U124 ( .A(n18), .B(n27), .Y(n278) );
  NAND2XL U125 ( .A(n108), .B(n11), .Y(n234) );
  NAND2XL U126 ( .A(a[7]), .B(n29), .Y(n450) );
  NAND2XL U127 ( .A(n100), .B(n104), .Y(n474) );
  NAND2XL U128 ( .A(n101), .B(n49), .Y(n222) );
  NAND2XL U129 ( .A(n18), .B(n102), .Y(n235) );
  NAND2XL U130 ( .A(n17), .B(n11), .Y(n303) );
  INVXL U131 ( .A(n107), .Y(n396) );
  NAND2XL U132 ( .A(n96), .B(n260), .Y(n263) );
  NOR2BXL U133 ( .AN(n111), .B(n30), .Y(n261) );
  XNOR3X2 U134 ( .A(n55), .B(n57), .C(n227), .Y(n228) );
  NAND2XL U135 ( .A(n36), .B(n18), .Y(n55) );
  NAND2XL U136 ( .A(n30), .B(n109), .Y(n57) );
  NAND2XL U137 ( .A(n101), .B(a[7]), .Y(n441) );
  NAND2XL U138 ( .A(n100), .B(a[7]), .Y(n401) );
  NAND2XL U139 ( .A(n100), .B(n47), .Y(n182) );
  NAND2XL U140 ( .A(a[5]), .B(n32), .Y(n499) );
  NAND2XL U141 ( .A(n101), .B(n23), .Y(n364) );
  NAND2XL U142 ( .A(n107), .B(n99), .Y(n363) );
  NAND2BXL U143 ( .AN(n100), .B(n110), .Y(n238) );
  NAND2XL U144 ( .A(a[3]), .B(n97), .Y(n482) );
  NAND2XL U145 ( .A(n105), .B(n98), .Y(n481) );
  XOR3X2 U146 ( .A(n58), .B(n416), .C(n375), .Y(n376) );
  NAND2XL U147 ( .A(a[1]), .B(n34), .Y(n58) );
  XOR3X2 U148 ( .A(n59), .B(n316), .C(n369), .Y(n317) );
  NAND2XL U149 ( .A(n31), .B(n26), .Y(n59) );
  XOR2X1 U150 ( .A(n60), .B(n61), .Y(n427) );
  XNOR3X2 U151 ( .A(n418), .B(n385), .C(n384), .Y(n60) );
  XNOR2X1 U152 ( .A(n420), .B(n419), .Y(n61) );
  NAND2XL U153 ( .A(n104), .B(n11), .Y(n428) );
  XOR3X2 U154 ( .A(n62), .B(n498), .C(n378), .Y(n339) );
  NAND2XL U155 ( .A(n104), .B(n30), .Y(n62) );
  XOR3X2 U156 ( .A(n63), .B(n362), .C(n361), .Y(n366) );
  NAND2XL U157 ( .A(n18), .B(b[2]), .Y(n63) );
  NAND2XL U158 ( .A(n11), .B(a[1]), .Y(n140) );
  NAND2XL U159 ( .A(n102), .B(a[3]), .Y(n142) );
  NAND2XL U160 ( .A(n100), .B(n17), .Y(n87) );
  NAND2XL U161 ( .A(n109), .B(n99), .Y(n92) );
  NAND2XL U162 ( .A(n17), .B(n99), .Y(n85) );
  NAND2XL U163 ( .A(n109), .B(n98), .Y(n86) );
  NAND2XL U164 ( .A(n30), .B(n26), .Y(n355) );
  NAND2BXL U165 ( .AN(b[2]), .B(n110), .Y(n148) );
  NAND2BXL U166 ( .AN(n30), .B(n33), .Y(n304) );
  NAND2BXL U167 ( .AN(n101), .B(n33), .Y(n260) );
  OAI2BB1X1 U168 ( .A0N(n110), .A1N(n119), .B0(n96), .Y(n126) );
  NAND2XL U169 ( .A(n106), .B(n11), .Y(n455) );
  NAND2XL U170 ( .A(n107), .B(n103), .Y(n456) );
  AND2X1 U171 ( .A(n47), .B(n98), .Y(n154) );
  AND2X1 U172 ( .A(n49), .B(n97), .Y(n139) );
  AND2X1 U173 ( .A(n109), .B(n102), .Y(n266) );
  XOR3X2 U174 ( .A(n64), .B(n410), .C(n95), .Y(n377) );
  NAND2XL U175 ( .A(a[3]), .B(n30), .Y(n64) );
  AND2X1 U176 ( .A(n31), .B(n105), .Y(n322) );
  AND2X1 U177 ( .A(n104), .B(n98), .Y(n219) );
  NAND2XL U178 ( .A(n12), .B(n105), .Y(n352) );
  NAND2XL U179 ( .A(a[5]), .B(n31), .Y(n371) );
  NAND2XL U180 ( .A(n31), .B(n23), .Y(n351) );
  NAND2XL U181 ( .A(a[4]), .B(n30), .Y(n431) );
  NAND2XL U182 ( .A(n23), .B(n37), .Y(n430) );
  NAND2XL U183 ( .A(b[4]), .B(a[5]), .Y(n507) );
  NAND2XL U184 ( .A(a[4]), .B(n31), .Y(n359) );
  NAND2XL U185 ( .A(n12), .B(n26), .Y(n319) );
  NAND2XL U186 ( .A(n23), .B(b[2]), .Y(n471) );
  NAND2XL U187 ( .A(n30), .B(n24), .Y(n360) );
  NAND2XL U188 ( .A(n13), .B(n23), .Y(n320) );
  NAND2XL U189 ( .A(a[4]), .B(n12), .Y(n370) );
  NAND2XL U190 ( .A(n24), .B(n34), .Y(n433) );
  NAND2XL U191 ( .A(b[1]), .B(n502), .Y(n65) );
  OAI2BB1X1 U192 ( .A0N(b[2]), .A1N(n136), .B0(n135), .Y(n138) );
  NAND2XL U193 ( .A(n96), .B(n133), .Y(n136) );
  NAND2BXL U194 ( .AN(b[1]), .B(n110), .Y(n133) );
  NAND2XL U195 ( .A(b[2]), .B(n49), .Y(n421) );
  AOI2BB2XL U196 ( .B0(b[0]), .B1(n387), .A0N(n96), .A1N(n501), .Y(n388) );
  NAND2XL U197 ( .A(b[0]), .B(n501), .Y(n66) );
  XNOR2X1 U198 ( .A(n147), .B(n179), .Y(n368) );
  XNOR2X1 U199 ( .A(n79), .B(n5), .Y(n321) );
  XOR2X1 U200 ( .A(n147), .B(n385), .Y(n67) );
  XOR3X2 U201 ( .A(n369), .B(n368), .C(n367), .Y(c[10]) );
  XOR2X1 U202 ( .A(n449), .B(n450), .Y(n178) );
  XNOR3X2 U203 ( .A(n67), .B(n180), .C(n213), .Y(n230) );
  XOR3X2 U204 ( .A(n214), .B(n290), .C(n213), .Y(n215) );
  XNOR3X2 U205 ( .A(n383), .B(n382), .C(n381), .Y(c[11]) );
  XNOR3X2 U206 ( .A(n372), .B(n371), .C(n370), .Y(n383) );
  XOR2X1 U207 ( .A(n377), .B(n376), .Y(n382) );
  XNOR3X2 U208 ( .A(n321), .B(n82), .C(n259), .Y(c[5]) );
  XNOR3X2 U209 ( .A(n470), .B(n254), .C(n253), .Y(n259) );
  XOR2X1 U210 ( .A(n252), .B(n471), .Y(n253) );
  XNOR2X1 U211 ( .A(n473), .B(n472), .Y(n254) );
  XNOR3X2 U212 ( .A(n347), .B(n346), .C(n343), .Y(c[8]) );
  XOR2X1 U213 ( .A(n320), .B(n319), .Y(n347) );
  XNOR2X1 U214 ( .A(n339), .B(n338), .Y(n343) );
  INVX1 U215 ( .A(n373), .Y(n385) );
  NOR2X1 U216 ( .A(n396), .B(n398), .Y(n418) );
  XOR3X2 U217 ( .A(n68), .B(n77), .C(n78), .Y(n367) );
  XNOR3X2 U218 ( .A(n409), .B(n408), .C(n407), .Y(n68) );
  XOR2X1 U219 ( .A(n360), .B(n359), .Y(n77) );
  XNOR2X1 U220 ( .A(n366), .B(n365), .Y(n78) );
  XOR2X1 U221 ( .A(n235), .B(n234), .Y(n251) );
  XOR3X2 U222 ( .A(n248), .B(n247), .C(n246), .Y(n249) );
  NAND2XL U223 ( .A(n202), .B(n196), .Y(n203) );
  INVX1 U224 ( .A(n375), .Y(n179) );
  XOR3X2 U225 ( .A(n80), .B(n81), .C(n228), .Y(n79) );
  XNOR2X1 U226 ( .A(n222), .B(n221), .Y(n80) );
  XOR2X1 U227 ( .A(n466), .B(n467), .Y(n81) );
  XOR2X1 U228 ( .A(n395), .B(n6), .Y(n378) );
  XNOR3X2 U229 ( .A(n83), .B(n296), .C(n292), .Y(c[6]) );
  XNOR3X2 U230 ( .A(n385), .B(n291), .C(n290), .Y(n292) );
  XOR2X1 U231 ( .A(n437), .B(n436), .Y(c[12]) );
  XOR2X1 U232 ( .A(n435), .B(n434), .Y(n436) );
  XOR2X1 U233 ( .A(n214), .B(n180), .Y(n82) );
  INVX1 U234 ( .A(n195), .Y(n196) );
  XNOR2X1 U235 ( .A(n301), .B(n5), .Y(n83) );
  XOR2X1 U236 ( .A(n318), .B(n317), .Y(c[7]) );
  XOR2X1 U237 ( .A(n216), .B(n215), .Y(c[3]) );
  XNOR3X2 U238 ( .A(n233), .B(n297), .C(n230), .Y(c[4]) );
  XNOR3X2 U239 ( .A(n83), .B(n358), .C(n357), .Y(c[9]) );
  NOR2XL U240 ( .A(n495), .B(n396), .Y(n488) );
  NAND4X1 U241 ( .A(n337), .B(n336), .C(n335), .D(n334), .Y(n395) );
  NAND3XL U242 ( .A(n37), .B(n331), .C(n333), .Y(n335) );
  OAI21XL U243 ( .A0(n15), .A1(n38), .B0(n50), .Y(n504) );
  OAI21XL U244 ( .A0(n18), .A1(n502), .B0(n66), .Y(n503) );
  OAI21XL U245 ( .A0(n23), .A1(n38), .B0(n50), .Y(n459) );
  OAI21XL U246 ( .A0(n105), .A1(n502), .B0(n7), .Y(n458) );
  XNOR2X1 U247 ( .A(n324), .B(n323), .Y(n333) );
  OAI21XL U248 ( .A0(n49), .A1(n38), .B0(n50), .Y(n405) );
  OAI21XL U249 ( .A0(n15), .A1(n502), .B0(n7), .Y(n406) );
  AOI22X1 U250 ( .A0(a[4]), .A1(n469), .B0(a[5]), .B1(n468), .Y(n470) );
  OAI21XL U251 ( .A0(n107), .A1(n38), .B0(n50), .Y(n469) );
  OAI21XL U252 ( .A0(n106), .A1(n502), .B0(n66), .Y(n468) );
  OAI21XL U253 ( .A0(n108), .A1(n501), .B0(n65), .Y(n478) );
  XNOR3X2 U254 ( .A(n453), .B(n454), .C(n210), .Y(n211) );
  NAND3X1 U255 ( .A(n205), .B(n204), .C(n203), .Y(n212) );
  NAND2X1 U256 ( .A(n20), .B(n37), .Y(n454) );
  OAI21XL U257 ( .A0(n107), .A1(n502), .B0(n7), .Y(n477) );
  OAI21XL U258 ( .A0(n26), .A1(n502), .B0(n66), .Y(n445) );
  OAI21XL U259 ( .A0(n23), .A1(n502), .B0(n66), .Y(n462) );
  OAI21XL U260 ( .A0(n21), .A1(n8), .B0(n7), .Y(n486) );
  XOR2X1 U261 ( .A(n166), .B(n165), .Y(n180) );
  XNOR3X2 U262 ( .A(n442), .B(n164), .C(n163), .Y(n165) );
  XNOR3X2 U263 ( .A(n154), .B(n153), .C(n152), .Y(n166) );
  INVX1 U264 ( .A(b[2]), .Y(n495) );
  XOR3X2 U265 ( .A(n188), .B(n187), .C(n182), .Y(n195) );
  NAND2X1 U266 ( .A(n29), .B(n17), .Y(n187) );
  NAND2X1 U267 ( .A(n101), .B(n109), .Y(n188) );
  XOR2X1 U268 ( .A(n289), .B(n288), .Y(n301) );
  XOR2X1 U269 ( .A(n286), .B(n278), .Y(n288) );
  XNOR3X2 U270 ( .A(n266), .B(n265), .C(n264), .Y(n289) );
  OAI2BB1X1 U271 ( .A0N(n11), .A1N(n132), .B0(n131), .Y(n375) );
  OAI21XL U272 ( .A0(n130), .A1(n387), .B0(n27), .Y(n131) );
  OAI2BB1X1 U273 ( .A0N(n33), .A1N(n129), .B0(n386), .Y(n132) );
  NOR2BX1 U274 ( .AN(n14), .B(n11), .Y(n130) );
  NOR2BX1 U275 ( .AN(n110), .B(n97), .Y(n170) );
  XOR2X1 U276 ( .A(n146), .B(n145), .Y(n213) );
  XNOR3X2 U277 ( .A(n400), .B(n144), .C(n143), .Y(n145) );
  XNOR3X2 U278 ( .A(n139), .B(n138), .C(n137), .Y(n146) );
  XNOR3X2 U279 ( .A(n384), .B(n350), .C(n349), .Y(n358) );
  XOR2X1 U280 ( .A(n348), .B(n507), .Y(n349) );
  XNOR2X1 U281 ( .A(n508), .B(n505), .Y(n350) );
  NAND2X1 U282 ( .A(a[4]), .B(n13), .Y(n348) );
  NAND2X1 U283 ( .A(b[4]), .B(n20), .Y(n416) );
  XOR2X1 U284 ( .A(n300), .B(n299), .Y(n316) );
  NAND2X1 U285 ( .A(n104), .B(n12), .Y(n299) );
  AND2X2 U286 ( .A(n106), .B(n103), .Y(n84) );
  XOR2X1 U287 ( .A(n169), .B(n168), .Y(n176) );
  XOR2X1 U288 ( .A(n162), .B(n155), .Y(n164) );
  XOR2X1 U289 ( .A(n402), .B(n403), .Y(n144) );
  NAND2X1 U290 ( .A(n106), .B(n36), .Y(n402) );
  XOR3X2 U291 ( .A(n428), .B(n429), .C(n395), .Y(n437) );
  XOR2X1 U292 ( .A(n425), .B(n424), .Y(n426) );
  XNOR3X2 U293 ( .A(n489), .B(n298), .C(n297), .Y(n318) );
  XOR3X2 U294 ( .A(n490), .B(n491), .C(n488), .Y(n298) );
  AOI22X1 U295 ( .A0(n21), .A1(n487), .B0(n20), .B1(n486), .Y(n489) );
  NAND2X1 U296 ( .A(n106), .B(n32), .Y(n491) );
  XNOR3X2 U297 ( .A(n67), .B(n457), .C(n181), .Y(n216) );
  NOR2X1 U298 ( .A(n397), .B(n399), .Y(n457) );
  XNOR2X1 U299 ( .A(n460), .B(n461), .Y(n181) );
  INVX1 U300 ( .A(n97), .Y(n399) );
  XOR2X1 U301 ( .A(n423), .B(n422), .Y(n424) );
  XOR2X1 U302 ( .A(n482), .B(n481), .Y(n483) );
  NAND2X1 U303 ( .A(n106), .B(b[4]), .Y(n498) );
  OAI2BB1X1 U304 ( .A0N(n110), .A1N(n223), .B0(n96), .Y(n226) );
  NAND2X1 U305 ( .A(n108), .B(n36), .Y(n449) );
  NAND2X1 U306 ( .A(a[7]), .B(n27), .Y(n246) );
  NAND2X1 U307 ( .A(n108), .B(n103), .Y(n466) );
  OAI2BB1X1 U308 ( .A0N(n37), .A1N(n314), .B0(n306), .Y(n315) );
  OAI21XL U309 ( .A0(n305), .A1(n387), .B0(n30), .Y(n306) );
  NOR2BX1 U310 ( .AN(n14), .B(n37), .Y(n305) );
  OAI2BB1X1 U311 ( .A0N(n97), .A1N(n174), .B0(n173), .Y(n175) );
  OAI21XL U312 ( .A0(n170), .A1(n189), .B0(n98), .Y(n173) );
  NAND2BX1 U313 ( .AN(n66), .B(n14), .Y(n389) );
  XNOR3X2 U314 ( .A(n85), .B(n86), .C(n401), .Y(n137) );
  XOR3X2 U315 ( .A(n142), .B(n141), .C(n140), .Y(n143) );
  NAND2X1 U316 ( .A(n103), .B(n105), .Y(n141) );
  XOR2X1 U317 ( .A(n448), .B(n447), .Y(n452) );
  NOR2X1 U318 ( .A(n397), .B(n495), .Y(n447) );
  AOI22X1 U319 ( .A0(n26), .A1(n446), .B0(n24), .B1(n445), .Y(n448) );
  OAI21XL U320 ( .A0(n105), .A1(n38), .B0(n50), .Y(n446) );
  XNOR3X2 U321 ( .A(n356), .B(n355), .C(n354), .Y(n357) );
  XOR3X2 U322 ( .A(n353), .B(n352), .C(n351), .Y(n354) );
  XOR2X1 U323 ( .A(n395), .B(n506), .Y(n356) );
  AOI21X1 U324 ( .A0(n100), .A1(n226), .B0(n225), .Y(n227) );
  OAI2BB1X1 U325 ( .A0N(n30), .A1N(n263), .B0(n262), .Y(n264) );
  OAI21XL U326 ( .A0(n261), .A1(n387), .B0(n101), .Y(n262) );
  XNOR3X2 U327 ( .A(n404), .B(n368), .C(n213), .Y(c[0]) );
  NOR2X1 U328 ( .A(n397), .B(n8), .Y(n404) );
  XOR2X1 U329 ( .A(n480), .B(n479), .Y(n484) );
  AOI22X1 U330 ( .A0(n107), .A1(n478), .B0(n108), .B1(n477), .Y(n480) );
  NAND2X1 U331 ( .A(n99), .B(n20), .Y(n420) );
  XOR2X1 U332 ( .A(n485), .B(n476), .Y(n296) );
  XOR2X1 U333 ( .A(n475), .B(n474), .Y(n476) );
  XOR2X1 U334 ( .A(n484), .B(n483), .Y(n485) );
  NAND2X1 U335 ( .A(n99), .B(a[1]), .Y(n475) );
  INVX1 U336 ( .A(n191), .Y(n194) );
  OAI21XL U337 ( .A0(n190), .A1(n189), .B0(n99), .Y(n191) );
  NOR2BX1 U338 ( .AN(n110), .B(n98), .Y(n190) );
  INVX1 U339 ( .A(n193), .Y(n202) );
  OAI21XL U340 ( .A0(n192), .A1(n387), .B0(n98), .Y(n193) );
  NOR2BX1 U341 ( .AN(n14), .B(n99), .Y(n192) );
  OAI21XL U342 ( .A0(n18), .A1(n38), .B0(n50), .Y(n493) );
  OAI21XL U343 ( .A0(n20), .A1(n502), .B0(n7), .Y(n492) );
  OAI21XL U344 ( .A0(n33), .A1(n38), .B0(n50), .Y(n412) );
  OAI21XL U345 ( .A0(n49), .A1(n8), .B0(n66), .Y(n411) );
  XOR2X1 U346 ( .A(n465), .B(n220), .Y(n233) );
  XOR3X2 U347 ( .A(n219), .B(n217), .C(n464), .Y(n220) );
  AOI22XL U348 ( .A0(n23), .A1(n463), .B0(n106), .B1(n462), .Y(n465) );
  NOR2X1 U349 ( .A(n495), .B(n500), .Y(n464) );
  INVX1 U350 ( .A(n102), .Y(n119) );
  NAND2BXL U351 ( .AN(n101), .B(n111), .Y(n237) );
  OAI2BB1X1 U352 ( .A0N(n97), .A1N(n151), .B0(n150), .Y(n153) );
  OAI21XL U353 ( .A0(n149), .A1(n387), .B0(b[2]), .Y(n150) );
  NOR2BX1 U354 ( .AN(n111), .B(n97), .Y(n149) );
  AND2X2 U355 ( .A(n10), .B(a[3]), .Y(n167) );
  XNOR3X2 U356 ( .A(n87), .B(n92), .C(n441), .Y(n152) );
  AND2X2 U357 ( .A(n47), .B(n99), .Y(n177) );
  XNOR2X1 U358 ( .A(n443), .B(n440), .Y(n163) );
  XNOR2X1 U359 ( .A(n455), .B(n456), .Y(n210) );
  INVX1 U360 ( .A(n99), .Y(n223) );
  INVX1 U361 ( .A(n103), .Y(n129) );
  OAI21XL U362 ( .A0(n106), .A1(n38), .B0(n50), .Y(n463) );
  OAI21XL U363 ( .A0(n20), .A1(n38), .B0(n50), .Y(n487) );
  NAND2X1 U364 ( .A(n105), .B(n37), .Y(n410) );
  XOR2X1 U365 ( .A(n374), .B(n373), .Y(n95) );
  NAND2X1 U366 ( .A(n104), .B(n34), .Y(n361) );
  NAND2X1 U367 ( .A(n37), .B(a[1]), .Y(n362) );
  XOR2X1 U368 ( .A(n364), .B(n363), .Y(n365) );
  XOR2X1 U369 ( .A(n433), .B(n432), .Y(n434) );
  NAND2X1 U370 ( .A(n26), .B(n27), .Y(n432) );
  XOR2X1 U371 ( .A(n499), .B(n496), .Y(n338) );
  NOR2X1 U372 ( .A(n495), .B(n494), .Y(n496) );
  INVX1 U373 ( .A(n108), .Y(n494) );
  AND2X2 U374 ( .A(n97), .B(a[1]), .Y(n217) );
  NAND2X1 U375 ( .A(n13), .B(n24), .Y(n300) );
  NAND2X1 U376 ( .A(n104), .B(n13), .Y(n252) );
  NAND2X1 U377 ( .A(n32), .B(n21), .Y(n508) );
  NAND2X1 U378 ( .A(n104), .B(n27), .Y(n374) );
  NAND2X1 U379 ( .A(n105), .B(n32), .Y(n473) );
  AND2X2 U380 ( .A(n20), .B(b[2]), .Y(n505) );
  NAND2X1 U381 ( .A(n97), .B(n20), .Y(n409) );
  NAND2X1 U382 ( .A(n104), .B(n37), .Y(n353) );
  NAND2X1 U383 ( .A(n21), .B(n99), .Y(n372) );
  INVX1 U384 ( .A(n104), .Y(n397) );
  XOR2X1 U385 ( .A(n431), .B(n430), .Y(n435) );
  AOI22X1 U386 ( .A0(a[0]), .A1(n439), .B0(n26), .B1(n438), .Y(n444) );
  OAI21XL U387 ( .A0(n26), .A1(n38), .B0(n50), .Y(n439) );
  OAI21XL U388 ( .A0(a[0]), .A1(n8), .B0(n7), .Y(n438) );
  XOR2X1 U389 ( .A(n417), .B(n414), .Y(n380) );
  NOR2X1 U390 ( .A(n413), .B(n495), .Y(n414) );
  INVX1 U391 ( .A(n105), .Y(n500) );
  INVX1 U392 ( .A(b[0]), .Y(n502) );
  INVX1 U393 ( .A(b[1]), .Y(n501) );
  BUFX3 U394 ( .A(a[4]), .Y(n106) );
  BUFX3 U395 ( .A(a[6]), .Y(n108) );
  BUFX3 U396 ( .A(a[2]), .Y(n105) );
  BUFX3 U397 ( .A(a[5]), .Y(n107) );
  BUFX3 U398 ( .A(b[11]), .Y(n103) );
  BUFX3 U399 ( .A(a[9]), .Y(n109) );
  BUFX3 U400 ( .A(b[10]), .Y(n102) );
  BUFX3 U401 ( .A(b[4]), .Y(n98) );
  BUFX3 U402 ( .A(b[7]), .Y(n101) );
  BUFX3 U403 ( .A(b[3]), .Y(n97) );
  BUFX3 U404 ( .A(b[5]), .Y(n99) );
  BUFX3 U405 ( .A(b[6]), .Y(n100) );
  XOR2X1 U406 ( .A(n394), .B(n421), .Y(n425) );
  OAI21XL U407 ( .A0(n134), .A1(n387), .B0(b[1]), .Y(n135) );
  NOR2BX1 U408 ( .AN(n111), .B(b[2]), .Y(n134) );
  BUFX3 U409 ( .A(a[0]), .Y(n104) );
  NAND2XL U410 ( .A(n327), .B(n326), .Y(n331) );
  AOI21XL U411 ( .A0(n327), .A1(n237), .B0(n236), .Y(n240) );
  AOI21XL U412 ( .A0(n327), .A1(n224), .B0(n223), .Y(n225) );
endmodule


module multiplier_8 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n36, n37, n38, n39, n47, n49, n50, n51, n52, n53,
         n54, n55, n57, n58, n59, n61, n63, n64, n74, n77, n81, n83, n84, n85,
         n86, n87, n92, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n122, n127, n128, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n202, n203, n204, n205, n210,
         n211, n212, n213, n214, n215, n216, n217, n219, n220, n221, n239,
         n240, n246, n247, n248, n249, n250, n251, n252, n253, n254, n259,
         n260, n261, n262, n263, n264, n265, n266, n286, n288, n289, n290,
         n291, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n311, n314, n315, n316, n317, n318, n319, n320, n321, n323,
         n324, n325, n326, n327, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540;

  CLKINVX3 U1 ( .A(n212), .Y(n217) );
  INVX1 U2 ( .A(n138), .Y(n332) );
  OAI21XL U3 ( .A0(n376), .A1(n375), .B0(n374), .Y(n450) );
  AOI21X2 U4 ( .A0(n34), .A1(n103), .B0(n102), .Y(n104) );
  NOR2X1 U5 ( .A(n373), .B(n84), .Y(n164) );
  NOR2X1 U6 ( .A(n27), .B(n373), .Y(n220) );
  OAI2BB1X1 U7 ( .A0N(n26), .A1N(n37), .B0(n368), .Y(n303) );
  NOR2X1 U8 ( .A(n373), .B(n83), .Y(n128) );
  NOR2X1 U9 ( .A(n25), .B(n373), .Y(n301) );
  OAI2BB1X1 U10 ( .A0N(n36), .A1N(n316), .B0(n368), .Y(n103) );
  AND2X2 U11 ( .A(n83), .B(n100), .Y(n521) );
  NOR2X1 U12 ( .A(n168), .B(n169), .Y(n1) );
  INVX1 U13 ( .A(n1), .Y(n170) );
  OAI221XL U14 ( .A0(n105), .A1(n58), .B0(n2), .B1(n373), .C0(n369), .Y(n370)
         );
  NOR2X1 U15 ( .A(n520), .B(n13), .Y(n413) );
  XNOR2X1 U16 ( .A(n380), .B(n215), .Y(n362) );
  OR2X2 U17 ( .A(n169), .B(n165), .Y(n174) );
  XNOR2X1 U18 ( .A(n138), .B(n215), .Y(n366) );
  OAI21XL U19 ( .A0(n375), .A1(n140), .B0(n83), .Y(n141) );
  INVX1 U20 ( .A(n315), .Y(n375) );
  NAND3X1 U21 ( .A(n169), .B(n165), .C(n168), .Y(n173) );
  OAI21XL U22 ( .A0(b[10]), .A1(n373), .B0(n315), .Y(n319) );
  XOR3X2 U23 ( .A(n352), .B(n336), .C(n351), .Y(c[10]) );
  XNOR3X2 U24 ( .A(n378), .B(n467), .C(n180), .Y(c[2]) );
  NOR2X1 U25 ( .A(n371), .B(n394), .Y(n372) );
  INVX1 U26 ( .A(b[3]), .Y(n394) );
  XOR2X1 U27 ( .A(n466), .B(n465), .Y(n494) );
  INVX1 U28 ( .A(n494), .Y(n383) );
  AOI21XL U29 ( .A0(n315), .A1(n259), .B0(n254), .Y(n262) );
  XOR2X4 U30 ( .A(n104), .B(n77), .Y(n138) );
  NAND2BX1 U31 ( .AN(a[11]), .B(a[12]), .Y(n315) );
  NAND2BX1 U32 ( .AN(a[12]), .B(n36), .Y(n166) );
  INVX1 U33 ( .A(n373), .Y(n32) );
  BUFX3 U34 ( .A(a[11]), .Y(n36) );
  BUFX3 U35 ( .A(n368), .Y(n81) );
  INVX1 U36 ( .A(a[12]), .Y(n373) );
  NAND2X1 U37 ( .A(b[0]), .B(n532), .Y(n2) );
  NAND2X1 U38 ( .A(b[0]), .B(n532), .Y(n57) );
  BUFX3 U39 ( .A(n58), .Y(n3) );
  NAND2X1 U40 ( .A(b[1]), .B(n533), .Y(n58) );
  INVX1 U41 ( .A(b[0]), .Y(n4) );
  INVX1 U42 ( .A(n389), .Y(n5) );
  BUFX3 U43 ( .A(b[3]), .Y(n6) );
  INVX1 U44 ( .A(n385), .Y(n7) );
  INVX1 U45 ( .A(n388), .Y(n8) );
  INVX1 U46 ( .A(n190), .Y(n9) );
  INVX1 U47 ( .A(a[10]), .Y(n10) );
  INVX1 U48 ( .A(n10), .Y(n11) );
  INVX1 U49 ( .A(n10), .Y(n12) );
  INVX1 U50 ( .A(a[9]), .Y(n13) );
  INVX1 U51 ( .A(n13), .Y(n14) );
  INVX1 U52 ( .A(n13), .Y(n15) );
  INVX1 U53 ( .A(a[8]), .Y(n16) );
  INVX1 U54 ( .A(n16), .Y(n17) );
  INVX1 U55 ( .A(n16), .Y(n18) );
  INVX1 U56 ( .A(a[7]), .Y(n19) );
  INVXL U57 ( .A(n19), .Y(n20) );
  INVX1 U58 ( .A(n500), .Y(n21) );
  INVX1 U59 ( .A(n531), .Y(n22) );
  INVX1 U60 ( .A(b[9]), .Y(n23) );
  INVX1 U61 ( .A(n23), .Y(n24) );
  INVX1 U62 ( .A(n23), .Y(n25) );
  INVX1 U63 ( .A(b[8]), .Y(n26) );
  INVX1 U64 ( .A(n26), .Y(n27) );
  INVXL U65 ( .A(n26), .Y(n28) );
  INVX1 U66 ( .A(n254), .Y(n29) );
  OAI21XL U67 ( .A0(n100), .A1(n367), .B0(n58), .Y(n499) );
  XOR2X4 U68 ( .A(n151), .B(n150), .Y(n378) );
  XNOR3X4 U69 ( .A(n145), .B(n144), .C(n143), .Y(n151) );
  BUFX3 U70 ( .A(b[10]), .Y(n30) );
  NAND2XL U71 ( .A(n18), .B(n30), .Y(n263) );
  INVX1 U72 ( .A(n464), .Y(n31) );
  NAND2XL U73 ( .A(n31), .B(n83), .Y(n487) );
  AOI22XL U74 ( .A0(n96), .A1(n474), .B0(n97), .B1(n473), .Y(n476) );
  NAND2X1 U75 ( .A(n97), .B(b[11]), .Y(n146) );
  NAND2BXL U76 ( .AN(n86), .B(n32), .Y(n259) );
  NOR2BXL U77 ( .AN(a[12]), .B(b[3]), .Y(n140) );
  NAND2BX1 U78 ( .AN(a[12]), .B(n37), .Y(n368) );
  BUFX3 U79 ( .A(b[4]), .Y(n33) );
  BUFX3 U80 ( .A(b[11]), .Y(n34) );
  CLKBUFX2 U81 ( .A(a[11]), .Y(n37) );
  XOR2X1 U82 ( .A(n493), .B(n492), .Y(c[5]) );
  XNOR3X2 U83 ( .A(n365), .B(n364), .C(n363), .Y(c[11]) );
  NAND2X1 U84 ( .A(n11), .B(n87), .Y(n77) );
  INVX1 U85 ( .A(n84), .Y(n190) );
  NAND2X1 U86 ( .A(n86), .B(n14), .Y(n163) );
  NAND2X1 U87 ( .A(n27), .B(n17), .Y(n162) );
  NAND2XL U88 ( .A(n97), .B(n6), .Y(n504) );
  NAND2XL U89 ( .A(n6), .B(n18), .Y(n416) );
  NAND2XL U90 ( .A(n98), .B(n6), .Y(n513) );
  NAND2XL U91 ( .A(n17), .B(n84), .Y(n61) );
  NAND2XL U92 ( .A(n6), .B(a[6]), .Y(n539) );
  AND2X1 U93 ( .A(n18), .B(n83), .Y(n404) );
  INVXL U94 ( .A(n366), .Y(n179) );
  XOR3X2 U95 ( .A(n39), .B(n286), .C(n266), .Y(n38) );
  XNOR2X1 U96 ( .A(n253), .B(n252), .Y(n39) );
  NOR2XL U97 ( .A(n385), .B(n389), .Y(n417) );
  NOR2XL U98 ( .A(n387), .B(n394), .Y(n472) );
  NOR2XL U99 ( .A(n386), .B(n389), .Y(n514) );
  XOR3X2 U100 ( .A(n47), .B(n404), .C(n49), .Y(n351) );
  XOR3X2 U101 ( .A(n405), .B(n338), .C(n337), .Y(n47) );
  XNOR3X2 U102 ( .A(n350), .B(n349), .C(n348), .Y(n49) );
  XOR2X1 U103 ( .A(n152), .B(n445), .Y(c[1]) );
  INVXL U104 ( .A(n36), .Y(n105) );
  AOI22XL U105 ( .A0(n8), .A1(n107), .B0(n34), .B1(n106), .Y(n380) );
  NAND2BXL U106 ( .AN(b[11]), .B(a[12]), .Y(n101) );
  NAND2XL U107 ( .A(n86), .B(n100), .Y(n397) );
  NAND2XL U108 ( .A(n25), .B(n11), .Y(n246) );
  NAND2XL U109 ( .A(n5), .B(n97), .Y(n338) );
  NAND2XL U110 ( .A(n86), .B(n18), .Y(n452) );
  AOI22XL U111 ( .A0(n18), .A1(n535), .B0(n15), .B1(n534), .Y(n537) );
  NAND2XL U112 ( .A(n98), .B(n24), .Y(n399) );
  NAND2XL U113 ( .A(n99), .B(n27), .Y(n400) );
  OAI21XL U114 ( .A0(n317), .A1(n371), .B0(n30), .Y(n318) );
  NAND2BXL U115 ( .AN(n85), .B(n32), .Y(n191) );
  INVXL U116 ( .A(n86), .Y(n389) );
  NAND2XL U117 ( .A(n20), .B(n8), .Y(n249) );
  NAND2XL U118 ( .A(n32), .B(n87), .Y(n215) );
  NAND2XL U119 ( .A(a[7]), .B(n25), .Y(n469) );
  OAI2BB1X1 U120 ( .A0N(b[3]), .A1N(n142), .B0(n141), .Y(n144) );
  NAND2XL U121 ( .A(n81), .B(n139), .Y(n142) );
  NAND2BXL U122 ( .AN(n83), .B(n37), .Y(n139) );
  NAND2XL U123 ( .A(b[4]), .B(n20), .Y(n415) );
  NAND2XL U124 ( .A(n85), .B(n17), .Y(n64) );
  NAND2XL U125 ( .A(n14), .B(n84), .Y(n74) );
  NAND2XL U126 ( .A(n97), .B(b[4]), .Y(n512) );
  NAND2XL U127 ( .A(n33), .B(n99), .Y(n538) );
  XNOR3X2 U128 ( .A(n333), .B(n332), .C(n537), .Y(n334) );
  NAND2XL U129 ( .A(n83), .B(n12), .Y(n421) );
  NAND2XL U130 ( .A(n92), .B(n25), .Y(n330) );
  NAND2XL U131 ( .A(n86), .B(n96), .Y(n327) );
  NAND2XL U132 ( .A(n12), .B(n6), .Y(n135) );
  NAND2XL U133 ( .A(n85), .B(n100), .Y(n418) );
  NAND2XL U134 ( .A(n33), .B(n18), .Y(n422) );
  NAND2XL U135 ( .A(n98), .B(n33), .Y(n523) );
  NAND2XL U136 ( .A(n100), .B(n24), .Y(n456) );
  NAND2XL U137 ( .A(n28), .B(n95), .Y(n321) );
  NAND2XL U138 ( .A(n100), .B(n34), .Y(n482) );
  NAND2XL U139 ( .A(n92), .B(n5), .Y(n296) );
  NAND2XL U140 ( .A(n29), .B(n92), .Y(n495) );
  NAND2XL U141 ( .A(a[7]), .B(b[11]), .Y(n252) );
  NAND2XL U142 ( .A(n98), .B(n34), .Y(n458) );
  NAND2XL U143 ( .A(n18), .B(n34), .Y(n248) );
  XOR3X2 U144 ( .A(n211), .B(n210), .C(n50), .Y(n384) );
  XNOR2X1 U145 ( .A(n205), .B(n204), .Y(n50) );
  NAND2XL U146 ( .A(n84), .B(n12), .Y(n451) );
  NAND2XL U147 ( .A(n17), .B(n87), .Y(n300) );
  NAND2XL U148 ( .A(n15), .B(b[11]), .Y(n299) );
  NAND2XL U149 ( .A(n87), .B(n96), .Y(n147) );
  NAND2XL U150 ( .A(n84), .B(n95), .Y(n496) );
  NAND2XL U151 ( .A(a[7]), .B(n30), .Y(n483) );
  NAND2XL U152 ( .A(n81), .B(n219), .Y(n239) );
  NAND2BXL U153 ( .AN(n86), .B(n37), .Y(n219) );
  NAND2XL U154 ( .A(n98), .B(n29), .Y(n339) );
  NAND2XL U155 ( .A(n25), .B(n95), .Y(n347) );
  NAND2XL U156 ( .A(n85), .B(a[7]), .Y(n398) );
  NAND2XL U157 ( .A(n86), .B(n20), .Y(n442) );
  NAND2XL U158 ( .A(n6), .B(n20), .Y(n407) );
  NAND2XL U159 ( .A(b[4]), .B(a[6]), .Y(n406) );
  NAND2XL U160 ( .A(n7), .B(n9), .Y(n337) );
  NAND2XL U161 ( .A(n85), .B(n11), .Y(n153) );
  NAND2BXL U162 ( .AN(n85), .B(n36), .Y(n260) );
  NAND2XL U163 ( .A(n6), .B(n15), .Y(n423) );
  NAND2XL U164 ( .A(a[7]), .B(n28), .Y(n457) );
  NAND2XL U165 ( .A(n96), .B(b[4]), .Y(n503) );
  NAND2XL U166 ( .A(n31), .B(n9), .Y(n516) );
  NAND2XL U167 ( .A(n29), .B(n96), .Y(n515) );
  NAND2XL U168 ( .A(n86), .B(n11), .Y(n195) );
  NAND2XL U169 ( .A(n27), .B(n14), .Y(n194) );
  AOI22XL U170 ( .A0(n12), .A1(n412), .B0(n36), .B1(n411), .Y(n414) );
  NAND2XL U171 ( .A(n85), .B(n97), .Y(n323) );
  XNOR3X2 U172 ( .A(n380), .B(n51), .C(n378), .Y(n381) );
  NAND2XL U173 ( .A(n84), .B(n92), .Y(n51) );
  XOR3X2 U174 ( .A(n52), .B(n306), .C(n336), .Y(n311) );
  NAND2XL U175 ( .A(n29), .B(a[1]), .Y(n52) );
  AOI22XL U176 ( .A0(a[6]), .A1(n509), .B0(n20), .B1(n508), .Y(n511) );
  NAND2XL U177 ( .A(n87), .B(n95), .Y(n108) );
  NAND2XL U178 ( .A(b[11]), .B(n96), .Y(n109) );
  NAND2XL U179 ( .A(n14), .B(n33), .Y(n63) );
  AOI22XL U180 ( .A0(n20), .A1(n519), .B0(n18), .B1(n518), .Y(n522) );
  NAND2XL U181 ( .A(n84), .B(n20), .Y(n419) );
  NAND2XL U182 ( .A(n92), .B(n8), .Y(n428) );
  NAND2XL U183 ( .A(n34), .B(n12), .Y(n410) );
  NAND2XL U184 ( .A(n98), .B(n87), .Y(n470) );
  NAND2XL U185 ( .A(n99), .B(n34), .Y(n471) );
  NAND2XL U186 ( .A(n99), .B(n24), .Y(n444) );
  NAND2XL U187 ( .A(n100), .B(n28), .Y(n441) );
  INVXL U188 ( .A(n87), .Y(n388) );
  INVX1 U189 ( .A(b[10]), .Y(n316) );
  AND2X1 U190 ( .A(n12), .B(n33), .Y(n145) );
  XNOR3X2 U191 ( .A(n53), .B(n410), .C(n320), .Y(n540) );
  NAND2XL U192 ( .A(n15), .B(n8), .Y(n53) );
  AND2X1 U193 ( .A(n14), .B(b[10]), .Y(n247) );
  AND2X1 U194 ( .A(n92), .B(b[4]), .Y(n188) );
  AND2X1 U195 ( .A(n98), .B(n84), .Y(n324) );
  XOR3X2 U196 ( .A(n55), .B(n305), .C(n304), .Y(n54) );
  NAND2XL U197 ( .A(n12), .B(n30), .Y(n55) );
  AND2X1 U198 ( .A(n20), .B(n83), .Y(n536) );
  INVX1 U199 ( .A(n166), .Y(n371) );
  XOR2X1 U200 ( .A(n455), .B(n454), .Y(n463) );
  XOR2X1 U201 ( .A(n453), .B(n452), .Y(n454) );
  NAND2XL U202 ( .A(n85), .B(n15), .Y(n453) );
  NAND2XL U203 ( .A(n99), .B(n87), .Y(n203) );
  NAND2XL U204 ( .A(n24), .B(n17), .Y(n202) );
  NAND2XL U205 ( .A(n28), .B(n96), .Y(n349) );
  NAND2XL U206 ( .A(n92), .B(n34), .Y(n359) );
  NAND2XL U207 ( .A(a[6]), .B(n9), .Y(n355) );
  NAND2XL U208 ( .A(n7), .B(n29), .Y(n356) );
  NAND2XL U209 ( .A(n21), .B(n5), .Y(n357) );
  NAND2XL U210 ( .A(n31), .B(n25), .Y(n431) );
  NAND2XL U211 ( .A(n31), .B(n28), .Y(n409) );
  NAND2XL U212 ( .A(n33), .B(n95), .Y(n488) );
  NAND2XL U213 ( .A(n95), .B(n34), .Y(n433) );
  NAND2XL U214 ( .A(n22), .B(n25), .Y(n408) );
  AND2X1 U215 ( .A(n28), .B(a[0]), .Y(n529) );
  NAND2XL U216 ( .A(n99), .B(n6), .Y(n524) );
  NAND2XL U217 ( .A(n22), .B(n30), .Y(n434) );
  NAND2XL U218 ( .A(a[1]), .B(n30), .Y(n358) );
  NAND2XL U219 ( .A(n21), .B(n28), .Y(n432) );
  NAND2XL U220 ( .A(n81), .B(n127), .Y(n132) );
  NAND2BXL U221 ( .AN(b[1]), .B(n37), .Y(n127) );
  AOI2BB2XL U222 ( .B0(b[0]), .B1(n375), .A0N(n81), .A1N(n367), .Y(n369) );
  INVXL U223 ( .A(b[1]), .Y(n367) );
  XOR2X1 U224 ( .A(n59), .B(n383), .Y(n288) );
  INVX1 U225 ( .A(n213), .Y(n152) );
  XOR2X1 U226 ( .A(n540), .B(n54), .Y(n354) );
  XOR2X1 U227 ( .A(n212), .B(n377), .Y(n290) );
  XNOR3X2 U228 ( .A(n179), .B(n178), .C(n378), .Y(n213) );
  XOR3X2 U229 ( .A(n265), .B(n264), .C(n263), .Y(n266) );
  XNOR3X2 U230 ( .A(n179), .B(n217), .C(n178), .Y(n181) );
  XOR2X1 U231 ( .A(n298), .B(n54), .Y(n336) );
  XNOR2X1 U232 ( .A(n494), .B(n380), .Y(n180) );
  XOR3X2 U233 ( .A(n514), .B(n38), .C(n384), .Y(n395) );
  XNOR3X2 U234 ( .A(n217), .B(n507), .C(n216), .Y(n289) );
  XOR2X1 U235 ( .A(n215), .B(n497), .Y(n216) );
  XOR2X1 U236 ( .A(n506), .B(n505), .Y(n507) );
  XOR2X1 U237 ( .A(n496), .B(n495), .Y(n497) );
  XOR3X2 U238 ( .A(n362), .B(n361), .C(n360), .Y(n363) );
  XOR2X1 U239 ( .A(n408), .B(n409), .Y(n361) );
  XNOR3X2 U240 ( .A(n415), .B(n359), .C(n358), .Y(n360) );
  INVX1 U241 ( .A(n384), .Y(n377) );
  XOR2X1 U242 ( .A(n289), .B(n288), .Y(c[6]) );
  XOR2X1 U243 ( .A(n438), .B(n437), .Y(c[12]) );
  XNOR2X1 U244 ( .A(n298), .B(n38), .Y(n59) );
  XOR2X1 U245 ( .A(n528), .B(n527), .Y(n530) );
  XOR2X1 U246 ( .A(n526), .B(n525), .Y(n527) );
  XOR2X1 U247 ( .A(n395), .B(n517), .Y(n528) );
  XOR2X1 U248 ( .A(n524), .B(n523), .Y(n525) );
  XOR2X1 U249 ( .A(n477), .B(n472), .Y(n182) );
  XOR2X1 U250 ( .A(n476), .B(n475), .Y(n477) );
  NOR2X1 U251 ( .A(n386), .B(n520), .Y(n475) );
  XOR3X2 U252 ( .A(n354), .B(n529), .C(n530), .Y(c[8]) );
  XOR2X1 U253 ( .A(n314), .B(n311), .Y(c[7]) );
  XNOR3X2 U254 ( .A(n182), .B(n181), .C(n180), .Y(c[3]) );
  XNOR3X2 U255 ( .A(n214), .B(n290), .C(n213), .Y(c[4]) );
  XNOR3X2 U256 ( .A(n335), .B(n59), .C(n334), .Y(c[9]) );
  NOR2X1 U257 ( .A(n520), .B(n385), .Y(n510) );
  OAI21XL U258 ( .A0(n34), .A1(n105), .B0(n81), .Y(n107) );
  OAI21XL U259 ( .A0(n15), .A1(n532), .B0(n3), .Y(n535) );
  OAI21XL U260 ( .A0(n18), .A1(n4), .B0(n57), .Y(n534) );
  OAI2BB1X1 U261 ( .A0N(n37), .A1N(n33), .B0(n394), .Y(n374) );
  MXI2X1 U262 ( .A(n373), .B(n372), .S0(b[4]), .Y(n376) );
  OAI21XL U263 ( .A0(n97), .A1(n367), .B0(n58), .Y(n474) );
  OAI21XL U264 ( .A0(n96), .A1(n4), .B0(n57), .Y(n473) );
  AOI22X1 U265 ( .A0(n12), .A1(n403), .B0(n15), .B1(n402), .Y(n405) );
  OAI21XL U266 ( .A0(n12), .A1(n367), .B0(n58), .Y(n402) );
  OAI21XL U267 ( .A0(n15), .A1(n4), .B0(n57), .Y(n403) );
  NOR2X1 U268 ( .A(n262), .B(n261), .Y(n286) );
  AOI21X1 U269 ( .A0(n81), .A1(n260), .B0(n389), .Y(n261) );
  INVXL U270 ( .A(n85), .Y(n254) );
  OAI2BB1X1 U271 ( .A0N(n25), .A1N(n319), .B0(n318), .Y(n320) );
  OAI21XL U272 ( .A0(n18), .A1(n367), .B0(n58), .Y(n519) );
  OAI21XL U273 ( .A0(n21), .A1(n367), .B0(n3), .Y(n479) );
  OAI21XL U274 ( .A0(n20), .A1(n367), .B0(n3), .Y(n509) );
  OAI21XL U275 ( .A0(n37), .A1(n367), .B0(n58), .Y(n412) );
  OAI21XL U276 ( .A0(n99), .A1(n4), .B0(n57), .Y(n498) );
  OAI21XL U277 ( .A0(n20), .A1(n4), .B0(n2), .Y(n518) );
  OAI21XL U278 ( .A0(n95), .A1(n4), .B0(n2), .Y(n446) );
  OAI21XL U279 ( .A0(n97), .A1(n4), .B0(n57), .Y(n478) );
  AOI22X1 U280 ( .A0(n21), .A1(n485), .B0(n7), .B1(n484), .Y(n486) );
  OAI21XL U281 ( .A0(n7), .A1(n367), .B0(n3), .Y(n485) );
  OAI21XL U282 ( .A0(n98), .A1(n533), .B0(n57), .Y(n484) );
  OAI21XL U283 ( .A0(a[6]), .A1(n533), .B0(n2), .Y(n508) );
  OAI21XL U284 ( .A0(n12), .A1(n4), .B0(n2), .Y(n411) );
  INVX1 U285 ( .A(n83), .Y(n520) );
  XNOR3X2 U286 ( .A(n443), .B(n149), .C(n148), .Y(n150) );
  NAND2X1 U287 ( .A(n98), .B(n30), .Y(n443) );
  OAI21XL U288 ( .A0(n301), .A1(n375), .B0(n28), .Y(n302) );
  XOR2X1 U289 ( .A(n137), .B(n136), .Y(n178) );
  XNOR3X2 U290 ( .A(n397), .B(n122), .C(n111), .Y(n137) );
  XNOR3X2 U291 ( .A(n135), .B(n134), .C(n133), .Y(n136) );
  XOR3X2 U292 ( .A(n163), .B(n162), .C(n153), .Y(n169) );
  XNOR2X1 U293 ( .A(n483), .B(n482), .Y(n210) );
  AOI21X1 U294 ( .A0(n85), .A1(n193), .B0(n192), .Y(n211) );
  XOR2X1 U295 ( .A(n177), .B(n176), .Y(n212) );
  XNOR3X2 U296 ( .A(n468), .B(n469), .C(n175), .Y(n176) );
  NAND3X1 U297 ( .A(n174), .B(n173), .C(n170), .Y(n177) );
  XOR2X1 U298 ( .A(n251), .B(n250), .Y(n298) );
  XOR2X1 U299 ( .A(n249), .B(n248), .Y(n250) );
  XNOR3X2 U300 ( .A(n247), .B(n246), .C(n240), .Y(n251) );
  NOR2X1 U301 ( .A(n388), .B(n464), .Y(n465) );
  XOR2X1 U302 ( .A(n463), .B(n462), .Y(n466) );
  INVX1 U303 ( .A(n97), .Y(n464) );
  NAND2X1 U304 ( .A(n100), .B(n87), .Y(n264) );
  XNOR2X1 U305 ( .A(n195), .B(n194), .Y(n205) );
  XOR2X1 U306 ( .A(n504), .B(n503), .Y(n505) );
  XOR3X2 U307 ( .A(n381), .B(n382), .C(n383), .Y(n492) );
  XOR2X1 U308 ( .A(n377), .B(n38), .Y(n382) );
  XOR2X1 U309 ( .A(n297), .B(n296), .Y(n306) );
  NAND2X1 U310 ( .A(n9), .B(n22), .Y(n297) );
  OAI2BB1X1 U311 ( .A0N(n25), .A1N(n303), .B0(n302), .Y(n304) );
  XOR2X1 U312 ( .A(n449), .B(n448), .Y(n467) );
  NOR2X1 U313 ( .A(n387), .B(n520), .Y(n448) );
  AOI22X1 U314 ( .A0(n95), .A1(n447), .B0(n22), .B1(n446), .Y(n449) );
  OAI21XL U315 ( .A0(n96), .A1(n367), .B0(n3), .Y(n447) );
  XOR2X1 U316 ( .A(n300), .B(n299), .Y(n305) );
  XOR2X1 U317 ( .A(n399), .B(n400), .Y(n122) );
  XOR2X1 U318 ( .A(n147), .B(n146), .Y(n149) );
  XNOR3X2 U319 ( .A(n511), .B(n291), .C(n290), .Y(n314) );
  XOR3X2 U320 ( .A(n512), .B(n513), .C(n510), .Y(n291) );
  XOR2X1 U321 ( .A(n203), .B(n202), .Y(n204) );
  XOR2X1 U322 ( .A(n461), .B(n460), .Y(n462) );
  XOR2X1 U323 ( .A(n457), .B(n456), .Y(n461) );
  XOR2X1 U324 ( .A(n459), .B(n458), .Y(n460) );
  XOR2X1 U325 ( .A(n425), .B(n424), .Y(n426) );
  XOR2X1 U326 ( .A(n423), .B(n422), .Y(n424) );
  XOR2X1 U327 ( .A(n370), .B(n421), .Y(n425) );
  OAI2BB1X1 U328 ( .A0N(n36), .A1N(n190), .B0(n81), .Y(n193) );
  NAND2X1 U329 ( .A(n27), .B(n11), .Y(n253) );
  XNOR3X2 U330 ( .A(n414), .B(n354), .C(n353), .Y(n365) );
  XNOR2X1 U331 ( .A(n413), .B(n416), .Y(n353) );
  NAND2X1 U332 ( .A(n99), .B(n30), .Y(n459) );
  XNOR3X2 U333 ( .A(n326), .B(n325), .C(n540), .Y(n335) );
  XOR2X1 U334 ( .A(n323), .B(n321), .Y(n326) );
  XOR2X1 U335 ( .A(n536), .B(n324), .Y(n325) );
  XNOR3X2 U336 ( .A(n61), .B(n63), .C(n398), .Y(n133) );
  XNOR3X2 U337 ( .A(n64), .B(n74), .C(n442), .Y(n143) );
  XOR3X2 U338 ( .A(n538), .B(n539), .C(n331), .Y(n333) );
  XNOR3X2 U339 ( .A(n110), .B(n109), .C(n108), .Y(n111) );
  NAND2X1 U340 ( .A(b[10]), .B(n97), .Y(n110) );
  NAND2X1 U341 ( .A(n24), .B(n15), .Y(n265) );
  NAND2X1 U342 ( .A(n100), .B(n30), .Y(n468) );
  OAI2BB1X1 U343 ( .A0N(n28), .A1N(n239), .B0(n221), .Y(n240) );
  OAI21XL U344 ( .A0(n220), .A1(n375), .B0(n86), .Y(n221) );
  XNOR3X2 U345 ( .A(n401), .B(n352), .C(n178), .Y(c[0]) );
  XOR2X1 U346 ( .A(n502), .B(n501), .Y(n506) );
  NOR2X1 U347 ( .A(n520), .B(n500), .Y(n501) );
  AOI22X1 U348 ( .A0(n99), .A1(n499), .B0(n100), .B1(n498), .Y(n502) );
  INVX1 U349 ( .A(n98), .Y(n500) );
  XOR2X1 U350 ( .A(n522), .B(n521), .Y(n526) );
  XOR2X1 U351 ( .A(n430), .B(n429), .Y(n438) );
  XNOR2X1 U352 ( .A(n428), .B(n540), .Y(n429) );
  XOR2X1 U353 ( .A(n427), .B(n426), .Y(n430) );
  XOR2X1 U354 ( .A(n451), .B(n450), .Y(n455) );
  XOR2X1 U355 ( .A(n396), .B(n420), .Y(n427) );
  XOR2X1 U356 ( .A(n419), .B(n418), .Y(n420) );
  XOR2X1 U357 ( .A(n366), .B(n417), .Y(n396) );
  XOR2X1 U358 ( .A(n491), .B(n490), .Y(n493) );
  XOR2X1 U359 ( .A(n489), .B(n488), .Y(n490) );
  XOR2X1 U360 ( .A(n487), .B(n486), .Y(n491) );
  NAND2X1 U361 ( .A(n22), .B(n6), .Y(n489) );
  OAI21XL U362 ( .A0(n164), .A1(n375), .B0(n33), .Y(n165) );
  OAI21XL U363 ( .A0(n167), .A1(n371), .B0(n84), .Y(n168) );
  NOR2BX1 U364 ( .AN(n36), .B(n33), .Y(n167) );
  XOR2X1 U365 ( .A(n481), .B(n189), .Y(n214) );
  XOR3X2 U366 ( .A(n188), .B(n187), .C(n480), .Y(n189) );
  AOI22X1 U367 ( .A0(n31), .A1(n479), .B0(n21), .B1(n478), .Y(n481) );
  NOR2X1 U368 ( .A(n520), .B(n531), .Y(n480) );
  XNOR2X1 U369 ( .A(n470), .B(n471), .Y(n175) );
  XNOR2X1 U370 ( .A(n444), .B(n441), .Y(n148) );
  NOR2BX1 U371 ( .AN(n36), .B(n25), .Y(n317) );
  AOI22X1 U372 ( .A0(a[0]), .A1(n440), .B0(a[1]), .B1(n439), .Y(n445) );
  OAI21XL U373 ( .A0(a[1]), .A1(n532), .B0(n3), .Y(n440) );
  OAI21XL U374 ( .A0(n92), .A1(n4), .B0(n2), .Y(n439) );
  NOR2X1 U375 ( .A(n387), .B(n4), .Y(n401) );
  XOR2X1 U376 ( .A(n516), .B(n515), .Y(n517) );
  XOR2X1 U377 ( .A(n436), .B(n435), .Y(n437) );
  XOR2X1 U378 ( .A(n432), .B(n431), .Y(n436) );
  XOR2X1 U379 ( .A(n434), .B(n433), .Y(n435) );
  AND2X2 U380 ( .A(n6), .B(n95), .Y(n187) );
  XOR3X2 U381 ( .A(n347), .B(n346), .C(n339), .Y(n348) );
  NAND2X1 U382 ( .A(n92), .B(n30), .Y(n346) );
  XNOR3X2 U383 ( .A(n357), .B(n356), .C(n355), .Y(n364) );
  INVX1 U384 ( .A(n92), .Y(n387) );
  XOR2X1 U385 ( .A(n330), .B(n327), .Y(n331) );
  XOR2X1 U386 ( .A(n407), .B(n406), .Y(n350) );
  INVX1 U387 ( .A(n95), .Y(n386) );
  INVX1 U388 ( .A(n99), .Y(n385) );
  INVX1 U389 ( .A(n96), .Y(n531) );
  OAI2BB1X1 U390 ( .A0N(n83), .A1N(n132), .B0(n131), .Y(n134) );
  OAI21XL U391 ( .A0(n128), .A1(n375), .B0(b[1]), .Y(n131) );
  BUFX3 U392 ( .A(a[3]), .Y(n97) );
  BUFX3 U393 ( .A(a[6]), .Y(n100) );
  BUFX3 U394 ( .A(a[2]), .Y(n96) );
  BUFX3 U395 ( .A(a[4]), .Y(n98) );
  BUFX3 U396 ( .A(a[5]), .Y(n99) );
  BUFX3 U397 ( .A(b[6]), .Y(n85) );
  BUFX3 U398 ( .A(a[1]), .Y(n95) );
  BUFX3 U399 ( .A(b[12]), .Y(n87) );
  BUFX3 U400 ( .A(b[7]), .Y(n86) );
  BUFX3 U401 ( .A(b[5]), .Y(n84) );
  INVX1 U402 ( .A(b[0]), .Y(n533) );
  INVX1 U403 ( .A(b[1]), .Y(n532) );
  BUFX3 U404 ( .A(b[2]), .Y(n83) );
  BUFX3 U405 ( .A(a[0]), .Y(n92) );
  OAI21XL U406 ( .A0(n87), .A1(n373), .B0(n315), .Y(n106) );
  AOI21X1 U407 ( .A0(n315), .A1(n191), .B0(n190), .Y(n192) );
  AOI21X1 U408 ( .A0(n315), .A1(n101), .B0(n316), .Y(n102) );
  XOR2X1 U409 ( .A(n138), .B(n380), .Y(n352) );
endmodule


module multiplier_7 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n47, n49, n50, n51, n52,
         n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n74, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n92,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n122, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n202,
         n203, n204, n205, n210, n211, n212, n213, n214, n215, n216, n217,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n230,
         n233, n234, n235, n236, n237, n238, n239, n240, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n259, n260, n261, n262, n263,
         n264, n265, n266, n278, n286, n288, n289, n290, n291, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n311, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n343, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502;

  CLKINVX3 U1 ( .A(n315), .Y(n378) );
  XOR2X2 U2 ( .A(n196), .B(n169), .Y(n65) );
  XOR2X2 U3 ( .A(n105), .B(n104), .Y(n374) );
  XOR2X1 U4 ( .A(n262), .B(n168), .Y(n196) );
  OAI21XL U5 ( .A0(n378), .A1(n101), .B0(n92), .Y(n102) );
  NOR2X1 U6 ( .A(n33), .B(n11), .Y(n104) );
  OAI21XL U7 ( .A0(n1), .A1(n87), .B0(n377), .Y(n249) );
  INVX1 U8 ( .A(n37), .Y(n1) );
  AOI211X1 U9 ( .A0(n317), .A1(n32), .B0(n322), .C0(n7), .Y(n2) );
  INVX1 U10 ( .A(n2), .Y(n325) );
  INVXL U11 ( .A(n319), .Y(n7) );
  NOR2X1 U12 ( .A(n489), .B(n25), .Y(n454) );
  NOR2XL U13 ( .A(n319), .B(n25), .Y(n80) );
  NOR2BX1 U14 ( .AN(n37), .B(n55), .Y(n382) );
  AND2X2 U15 ( .A(n82), .B(n100), .Y(n490) );
  OAI21XL U16 ( .A0(n3), .A1(n321), .B0(n322), .Y(n323) );
  INVX1 U17 ( .A(n320), .Y(n3) );
  NAND3XL U18 ( .A(n182), .B(n178), .C(n180), .Y(n190) );
  XNOR2X1 U19 ( .A(n220), .B(n438), .Y(c[1]) );
  INVX1 U20 ( .A(n374), .Y(n137) );
  NAND2X1 U21 ( .A(n99), .B(n92), .Y(n445) );
  CLKINVX3 U22 ( .A(n11), .Y(n13) );
  NAND2BX2 U23 ( .AN(a[11]), .B(a[12]), .Y(n315) );
  XOR2X1 U24 ( .A(n150), .B(n149), .Y(n169) );
  OAI2BB1X1 U25 ( .A0N(n95), .A1N(n103), .B0(n102), .Y(n105) );
  XOR2X4 U26 ( .A(n194), .B(n193), .Y(n261) );
  XOR2X1 U27 ( .A(n261), .B(n62), .Y(n265) );
  AND2X2 U28 ( .A(n97), .B(n32), .Y(n4) );
  XNOR3X2 U29 ( .A(n237), .B(n236), .C(n235), .Y(n5) );
  XNOR3X2 U30 ( .A(n47), .B(n49), .C(n299), .Y(n6) );
  NAND2XL U31 ( .A(b[1]), .B(n496), .Y(n8) );
  BUFX3 U32 ( .A(n57), .Y(n9) );
  INVX1 U33 ( .A(b[1]), .Y(n495) );
  INVX1 U34 ( .A(b[0]), .Y(n10) );
  INVX1 U35 ( .A(b[12]), .Y(n11) );
  INVX1 U36 ( .A(n11), .Y(n12) );
  INVX1 U37 ( .A(n387), .Y(n14) );
  INVX1 U38 ( .A(a[9]), .Y(n15) );
  INVX1 U39 ( .A(n15), .Y(n16) );
  INVX1 U40 ( .A(n15), .Y(n17) );
  INVX1 U41 ( .A(a[8]), .Y(n18) );
  INVX1 U42 ( .A(n18), .Y(n19) );
  INVX1 U43 ( .A(a[7]), .Y(n20) );
  INVXL U44 ( .A(n20), .Y(n21) );
  INVX1 U45 ( .A(a[3]), .Y(n22) );
  INVXL U46 ( .A(n22), .Y(n23) );
  INVX1 U47 ( .A(n494), .Y(n24) );
  INVX1 U48 ( .A(a[1]), .Y(n25) );
  INVX1 U49 ( .A(n25), .Y(n26) );
  INVX1 U50 ( .A(n106), .Y(n27) );
  INVX1 U51 ( .A(b[8]), .Y(n28) );
  INVX1 U52 ( .A(n28), .Y(n29) );
  INVX1 U53 ( .A(n224), .Y(n30) );
  INVX1 U54 ( .A(b[9]), .Y(n31) );
  INVX1 U55 ( .A(n31), .Y(n32) );
  AOI2BB2XL U56 ( .B0(b[0]), .B1(n378), .A0N(n81), .A1N(n376), .Y(n380) );
  NAND2BX1 U57 ( .AN(a[12]), .B(a[11]), .Y(n377) );
  BUFX3 U58 ( .A(n377), .Y(n81) );
  INVX1 U59 ( .A(a[10]), .Y(n33) );
  INVX1 U60 ( .A(n33), .Y(n34) );
  INVXL U61 ( .A(n33), .Y(n35) );
  BUFX3 U62 ( .A(a[12]), .Y(n36) );
  BUFX3 U63 ( .A(a[11]), .Y(n37) );
  OAI2BB1X2 U64 ( .A0N(a[11]), .A1N(n319), .B0(n81), .Y(n103) );
  NAND2X1 U65 ( .A(n34), .B(n95), .Y(n306) );
  NAND2X1 U66 ( .A(b[0]), .B(n495), .Y(n57) );
  XNOR3X2 U67 ( .A(n167), .B(n38), .C(n39), .Y(n262) );
  XNOR3X2 U68 ( .A(n151), .B(n445), .C(n68), .Y(n38) );
  XNOR3X2 U69 ( .A(n166), .B(n165), .C(n164), .Y(n39) );
  NOR2XL U70 ( .A(n54), .B(n319), .Y(n321) );
  INVXL U71 ( .A(n322), .Y(n318) );
  NAND2X1 U72 ( .A(n188), .B(n187), .Y(n189) );
  NAND2XL U73 ( .A(n187), .B(n181), .Y(n191) );
  XOR2X1 U74 ( .A(n65), .B(n446), .Y(c[2]) );
  INVXL U75 ( .A(n180), .Y(n188) );
  INVXL U76 ( .A(n95), .Y(n106) );
  OAI2BB1XL U77 ( .A0N(n37), .A1N(n106), .B0(n81), .Y(n109) );
  AOI22XL U78 ( .A0(n24), .A1(n453), .B0(n23), .B1(n452), .Y(n455) );
  AOI22XL U79 ( .A0(n19), .A1(n498), .B0(n17), .B1(n497), .Y(n500) );
  NAND2XL U80 ( .A(n87), .B(n100), .Y(n394) );
  AOI22XL U81 ( .A0(n35), .A1(n400), .B0(n17), .B1(n399), .Y(n401) );
  NAND2XL U82 ( .A(b[4]), .B(a[6]), .Y(n402) );
  NAND2XL U83 ( .A(n29), .B(n35), .Y(n233) );
  NAND2XL U84 ( .A(b[9]), .B(n35), .Y(n251) );
  NAND2BXL U85 ( .AN(n82), .B(a[11]), .Y(n138) );
  NAND2XL U86 ( .A(n81), .B(n138), .Y(n141) );
  NAND2BXL U87 ( .AN(n86), .B(n36), .Y(n214) );
  NAND2XL U88 ( .A(n35), .B(n92), .Y(n47) );
  XNOR2X1 U89 ( .A(n290), .B(n289), .Y(n49) );
  NAND2XL U90 ( .A(n12), .B(n97), .Y(n146) );
  NAND2XL U91 ( .A(a[3]), .B(n95), .Y(n145) );
  NAND2XL U92 ( .A(n98), .B(b[9]), .Y(n396) );
  NAND2XL U93 ( .A(n99), .B(b[8]), .Y(n397) );
  NAND2BXL U94 ( .AN(n92), .B(a[12]), .Y(n314) );
  NOR2X1 U95 ( .A(n228), .B(n227), .Y(n236) );
  AOI21XL U96 ( .A0(n81), .A1(n226), .B0(n387), .Y(n227) );
  NAND2XL U97 ( .A(a[7]), .B(n32), .Y(n448) );
  NAND2XL U98 ( .A(n36), .B(n13), .Y(n365) );
  NAND2XL U99 ( .A(n82), .B(n35), .Y(n415) );
  NAND2BXL U100 ( .AN(b[8]), .B(n37), .Y(n291) );
  NAND2XL U101 ( .A(n81), .B(n291), .Y(n298) );
  NAND2XL U102 ( .A(n21), .B(n27), .Y(n230) );
  NAND2XL U103 ( .A(n98), .B(n92), .Y(n436) );
  AOI22XL U104 ( .A0(n21), .A1(n488), .B0(n19), .B1(n487), .Y(n491) );
  NAND2XL U105 ( .A(n30), .B(n24), .Y(n67) );
  NAND2XL U106 ( .A(a[4]), .B(b[5]), .Y(n333) );
  NAND2XL U107 ( .A(n83), .B(n21), .Y(n403) );
  NAND2XL U108 ( .A(n100), .B(n92), .Y(n447) );
  NAND2XL U109 ( .A(a[3]), .B(n84), .Y(n485) );
  NAND2XL U110 ( .A(n86), .B(n34), .Y(n173) );
  NAND2XL U111 ( .A(b[8]), .B(a[8]), .Y(n174) );
  NAND2XL U112 ( .A(n87), .B(n16), .Y(n175) );
  NAND2XL U113 ( .A(b[9]), .B(n17), .Y(n234) );
  NAND2XL U114 ( .A(n32), .B(n317), .Y(n320) );
  NAND2XL U115 ( .A(n16), .B(n12), .Y(n311) );
  NAND2XL U116 ( .A(b[4]), .B(a[1]), .Y(n466) );
  INVXL U117 ( .A(n87), .Y(n387) );
  NAND2XL U118 ( .A(n99), .B(n13), .Y(n211) );
  NAND2XL U119 ( .A(n86), .B(n100), .Y(n412) );
  NAND2XL U120 ( .A(n100), .B(b[8]), .Y(n434) );
  NAND2XL U121 ( .A(n99), .B(b[9]), .Y(n437) );
  NAND2XL U122 ( .A(a[7]), .B(n7), .Y(n461) );
  NAND2XL U123 ( .A(n97), .B(n84), .Y(n476) );
  NAND2XL U124 ( .A(n16), .B(n95), .Y(n289) );
  NAND2XL U125 ( .A(n19), .B(n27), .Y(n253) );
  NAND2XL U126 ( .A(n100), .B(n13), .Y(n222) );
  NAND2XL U127 ( .A(a[7]), .B(b[8]), .Y(n444) );
  NOR2BXL U128 ( .AN(n36), .B(n13), .Y(n107) );
  NAND2XL U129 ( .A(b[3]), .B(a[6]), .Y(n502) );
  NAND2XL U130 ( .A(n87), .B(n35), .Y(n212) );
  NAND2XL U131 ( .A(n19), .B(n92), .Y(n223) );
  NAND2XL U132 ( .A(n97), .B(b[3]), .Y(n467) );
  NAND2XL U133 ( .A(n100), .B(n95), .Y(n460) );
  NAND2XL U134 ( .A(a[8]), .B(n12), .Y(n290) );
  AND2X1 U135 ( .A(n83), .B(a[1]), .Y(n204) );
  INVXL U136 ( .A(n99), .Y(n385) );
  NOR2BXL U137 ( .AN(a[11]), .B(n84), .Y(n177) );
  XNOR3X2 U138 ( .A(n50), .B(n51), .C(n217), .Y(n219) );
  NAND2XL U139 ( .A(n32), .B(n19), .Y(n50) );
  NAND2XL U140 ( .A(n29), .B(n17), .Y(n51) );
  NAND2XL U141 ( .A(n87), .B(a[7]), .Y(n435) );
  NAND2XL U142 ( .A(n86), .B(a[7]), .Y(n395) );
  NAND2BXL U143 ( .AN(n86), .B(n37), .Y(n226) );
  NAND2XL U144 ( .A(n87), .B(n23), .Y(n354) );
  NAND2XL U145 ( .A(n99), .B(n85), .Y(n353) );
  NAND2XL U146 ( .A(n83), .B(n17), .Y(n417) );
  NAND2XL U147 ( .A(n84), .B(n19), .Y(n416) );
  NAND2XL U148 ( .A(n85), .B(a[1]), .Y(n469) );
  NAND2XL U149 ( .A(n86), .B(n96), .Y(n468) );
  AOI22XL U150 ( .A0(n35), .A1(n406), .B0(n37), .B1(n405), .Y(n408) );
  NAND2XL U151 ( .A(b[3]), .B(n19), .Y(n410) );
  OAI2BB1XL U152 ( .A0N(n37), .A1N(n213), .B0(n81), .Y(n216) );
  XOR3X2 U153 ( .A(n52), .B(n300), .C(n359), .Y(n301) );
  NAND2XL U154 ( .A(n30), .B(n26), .Y(n52) );
  NAND2XL U155 ( .A(n96), .B(n13), .Y(n422) );
  AOI22XL U156 ( .A0(a[6]), .A1(n482), .B0(n21), .B1(n481), .Y(n484) );
  NAND2XL U157 ( .A(n98), .B(b[3]), .Y(n486) );
  INVXL U158 ( .A(n83), .Y(n388) );
  XOR3X2 U159 ( .A(n53), .B(n352), .C(n351), .Y(n356) );
  NAND2XL U160 ( .A(n19), .B(n82), .Y(n53) );
  NAND2XL U161 ( .A(n13), .B(a[1]), .Y(n130) );
  NAND2XL U162 ( .A(n95), .B(n97), .Y(n131) );
  NAND2XL U163 ( .A(n92), .B(a[3]), .Y(n132) );
  NAND2XL U164 ( .A(n86), .B(a[8]), .Y(n78) );
  NAND2XL U165 ( .A(n16), .B(n85), .Y(n79) );
  NAND2XL U166 ( .A(a[8]), .B(n85), .Y(n74) );
  NAND2XL U167 ( .A(n17), .B(n84), .Y(n77) );
  NAND2XL U168 ( .A(n29), .B(n26), .Y(n343) );
  NAND2XL U169 ( .A(a[3]), .B(n83), .Y(n477) );
  NAND2XL U170 ( .A(n85), .B(n21), .Y(n413) );
  XOR2X1 U171 ( .A(n260), .B(n259), .Y(n288) );
  NAND2XL U172 ( .A(n21), .B(n13), .Y(n254) );
  NAND2XL U173 ( .A(a[5]), .B(b[3]), .Y(n493) );
  NAND2XL U174 ( .A(n98), .B(n13), .Y(n449) );
  NAND2XL U175 ( .A(n99), .B(n95), .Y(n450) );
  NAND2XL U176 ( .A(n96), .B(n27), .Y(n366) );
  INVXL U177 ( .A(n85), .Y(n213) );
  AND2X1 U178 ( .A(n98), .B(n95), .Y(n68) );
  AND2X1 U179 ( .A(n34), .B(n84), .Y(n144) );
  AND2X1 U180 ( .A(n35), .B(n83), .Y(n129) );
  AND2X1 U181 ( .A(n17), .B(n92), .Y(n252) );
  AND2X1 U182 ( .A(n96), .B(n84), .Y(n205) );
  AND2X1 U183 ( .A(n96), .B(n29), .Y(n326) );
  AND2X1 U184 ( .A(n21), .B(n82), .Y(n499) );
  AND2X1 U185 ( .A(n81), .B(n316), .Y(n54) );
  NAND2XL U186 ( .A(n14), .B(n97), .Y(n337) );
  NAND2XL U187 ( .A(n98), .B(b[4]), .Y(n492) );
  NAND2XL U188 ( .A(n30), .B(n23), .Y(n336) );
  NAND2XL U189 ( .A(a[6]), .B(b[5]), .Y(n362) );
  NAND2XL U190 ( .A(a[5]), .B(n30), .Y(n363) );
  NAND2XL U191 ( .A(a[4]), .B(n14), .Y(n364) );
  NAND2XL U192 ( .A(b[4]), .B(n21), .Y(n409) );
  NAND2XL U193 ( .A(n96), .B(n32), .Y(n338) );
  NAND2XL U194 ( .A(n23), .B(n29), .Y(n404) );
  NAND2XL U195 ( .A(b[4]), .B(a[5]), .Y(n501) );
  NAND2XL U196 ( .A(n98), .B(n30), .Y(n349) );
  NAND2XL U197 ( .A(n96), .B(n14), .Y(n278) );
  NAND2XL U198 ( .A(n23), .B(n82), .Y(n465) );
  NAND2XL U199 ( .A(n29), .B(n97), .Y(n350) );
  NAND2XL U200 ( .A(a[0]), .B(b[5]), .Y(n238) );
  NAND2XL U201 ( .A(b[5]), .B(n23), .Y(n304) );
  NAND2XL U202 ( .A(n14), .B(n26), .Y(n303) );
  NAND2XL U203 ( .A(n24), .B(n7), .Y(n427) );
  NAND2XL U204 ( .A(n26), .B(n27), .Y(n426) );
  NAND2XL U205 ( .A(a[4]), .B(n29), .Y(n425) );
  NAND2XL U206 ( .A(n23), .B(n32), .Y(n424) );
  NAND2BXL U207 ( .AN(b[1]), .B(n37), .Y(n110) );
  NAND2XL U208 ( .A(n81), .B(n110), .Y(n126) );
  INVXL U209 ( .A(b[1]), .Y(n376) );
  NAND2X1 U210 ( .A(b[1]), .B(n496), .Y(n55) );
  XNOR2X1 U211 ( .A(n137), .B(n168), .Y(n358) );
  XNOR2X1 U212 ( .A(n62), .B(n5), .Y(n305) );
  XOR2X1 U213 ( .A(n137), .B(n375), .Y(n58) );
  XOR3X2 U214 ( .A(n359), .B(n358), .C(n357), .Y(c[10]) );
  NAND3X1 U215 ( .A(n325), .B(n324), .C(n323), .Y(n384) );
  NAND3X1 U216 ( .A(n54), .B(n318), .C(n320), .Y(n324) );
  XOR2X1 U217 ( .A(n443), .B(n444), .Y(n167) );
  XOR2X1 U218 ( .A(n384), .B(n6), .Y(n361) );
  XNOR3X2 U219 ( .A(n58), .B(n169), .C(n195), .Y(n220) );
  XNOR3X2 U220 ( .A(n332), .B(n331), .C(n330), .Y(c[8]) );
  XOR3X2 U221 ( .A(n196), .B(n261), .C(n195), .Y(n202) );
  XNOR3X2 U222 ( .A(n305), .B(n65), .C(n246), .Y(c[5]) );
  XNOR3X2 U223 ( .A(n464), .B(n240), .C(n239), .Y(n246) );
  XOR2X1 U224 ( .A(n238), .B(n465), .Y(n239) );
  XNOR2X1 U225 ( .A(n467), .B(n466), .Y(n240) );
  INVX1 U226 ( .A(n365), .Y(n375) );
  NOR2X1 U227 ( .A(n385), .B(n387), .Y(n411) );
  XNOR3X2 U228 ( .A(n221), .B(n265), .C(n220), .Y(c[4]) );
  XOR3X2 U229 ( .A(n59), .B(n60), .C(n61), .Y(n357) );
  XNOR3X2 U230 ( .A(n403), .B(n402), .C(n401), .Y(n59) );
  XOR2X1 U231 ( .A(n350), .B(n349), .Y(n60) );
  XNOR2X1 U232 ( .A(n356), .B(n355), .Y(n61) );
  INVX1 U233 ( .A(n368), .Y(n168) );
  XOR2X1 U234 ( .A(n223), .B(n222), .Y(n237) );
  XOR3X2 U235 ( .A(n234), .B(n233), .C(n230), .Y(n235) );
  XNOR3X2 U236 ( .A(n375), .B(n262), .C(n261), .Y(n263) );
  XOR3X2 U237 ( .A(n63), .B(n64), .C(n219), .Y(n62) );
  XNOR2X1 U238 ( .A(n212), .B(n211), .Y(n63) );
  XOR2X1 U239 ( .A(n460), .B(n461), .Y(n64) );
  XNOR3X2 U240 ( .A(n66), .B(n264), .C(n263), .Y(c[6]) );
  XOR2X1 U241 ( .A(n480), .B(n470), .Y(n264) );
  XOR2X1 U242 ( .A(n431), .B(n430), .Y(c[12]) );
  XOR2X1 U243 ( .A(n429), .B(n428), .Y(n430) );
  XOR2X1 U244 ( .A(n370), .B(n369), .Y(n371) );
  XNOR3X2 U245 ( .A(n404), .B(n4), .C(n367), .Y(n370) );
  XOR3X2 U246 ( .A(n409), .B(n368), .C(n80), .Y(n369) );
  INVX1 U247 ( .A(n182), .Y(n187) );
  INVX1 U248 ( .A(n377), .Y(n176) );
  XNOR2X1 U249 ( .A(n288), .B(n5), .Y(n66) );
  XOR2XL U250 ( .A(n288), .B(n6), .Y(n359) );
  XOR2X1 U251 ( .A(n302), .B(n301), .Y(c[7]) );
  XOR2X1 U252 ( .A(n203), .B(n202), .Y(c[3]) );
  XNOR3X2 U253 ( .A(n66), .B(n348), .C(n347), .Y(c[9]) );
  XOR3X2 U254 ( .A(n373), .B(n372), .C(n371), .Y(c[11]) );
  NOR2XL U255 ( .A(n489), .B(n385), .Y(n483) );
  OAI21XL U256 ( .A0(n17), .A1(n376), .B0(n8), .Y(n498) );
  OAI21XL U257 ( .A0(n19), .A1(n496), .B0(n57), .Y(n497) );
  OAI21XL U258 ( .A0(n23), .A1(n495), .B0(n8), .Y(n453) );
  OAI21XL U259 ( .A0(n97), .A1(n10), .B0(n57), .Y(n452) );
  AOI22X1 U260 ( .A0(n99), .A1(n472), .B0(n100), .B1(n471), .Y(n475) );
  OAI21XL U261 ( .A0(n100), .A1(n376), .B0(n55), .Y(n472) );
  OAI21XL U262 ( .A0(n99), .A1(n496), .B0(n57), .Y(n471) );
  OAI21XL U263 ( .A0(n35), .A1(n376), .B0(n8), .Y(n399) );
  OAI21XL U264 ( .A0(n17), .A1(n10), .B0(n57), .Y(n400) );
  OAI2BB1X1 U265 ( .A0N(n13), .A1N(n109), .B0(n108), .Y(n368) );
  INVXL U266 ( .A(n86), .Y(n224) );
  OAI21XL U267 ( .A0(n26), .A1(n10), .B0(n9), .Y(n439) );
  OAI21XL U268 ( .A0(n21), .A1(n10), .B0(n57), .Y(n487) );
  OAI21XL U269 ( .A0(n23), .A1(n10), .B0(n9), .Y(n456) );
  AOI22X1 U270 ( .A0(a[4]), .A1(n463), .B0(a[5]), .B1(n462), .Y(n464) );
  OAI21XL U271 ( .A0(n99), .A1(n376), .B0(n8), .Y(n463) );
  OAI21XL U272 ( .A0(n98), .A1(n10), .B0(n57), .Y(n462) );
  OAI21XL U273 ( .A0(a[6]), .A1(n10), .B0(n57), .Y(n481) );
  OAI21XL U274 ( .A0(n35), .A1(n10), .B0(n57), .Y(n405) );
  OAI21XL U275 ( .A0(n19), .A1(n376), .B0(n8), .Y(n488) );
  OAI21XL U276 ( .A0(n37), .A1(n376), .B0(n8), .Y(n406) );
  XNOR3X2 U277 ( .A(n436), .B(n148), .C(n147), .Y(n149) );
  XNOR3X2 U278 ( .A(n144), .B(n143), .C(n142), .Y(n150) );
  NOR2X1 U279 ( .A(n489), .B(n473), .Y(n474) );
  INVX1 U280 ( .A(n98), .Y(n473) );
  INVX1 U281 ( .A(n82), .Y(n489) );
  XNOR3X2 U282 ( .A(n447), .B(n448), .C(n192), .Y(n193) );
  NAND3X1 U283 ( .A(n191), .B(n190), .C(n189), .Y(n194) );
  OAI2BB1X1 U284 ( .A0N(n83), .A1N(n141), .B0(n140), .Y(n143) );
  XOR2X1 U285 ( .A(n254), .B(n253), .Y(n259) );
  XNOR3X2 U286 ( .A(n252), .B(n251), .C(n250), .Y(n260) );
  NOR2BX1 U287 ( .AN(a[12]), .B(n95), .Y(n101) );
  NOR2BX1 U288 ( .AN(a[11]), .B(n83), .Y(n155) );
  XNOR2X1 U289 ( .A(n311), .B(n306), .Y(n322) );
  XOR2X1 U290 ( .A(n136), .B(n135), .Y(n195) );
  XNOR3X2 U291 ( .A(n394), .B(n134), .C(n133), .Y(n135) );
  XNOR3X2 U292 ( .A(n129), .B(n128), .C(n127), .Y(n136) );
  XNOR3X2 U293 ( .A(n374), .B(n335), .C(n334), .Y(n348) );
  XOR2X1 U294 ( .A(n333), .B(n501), .Y(n334) );
  XNOR2X1 U295 ( .A(n502), .B(n499), .Y(n335) );
  XNOR3X2 U296 ( .A(n67), .B(n491), .C(n305), .Y(n331) );
  NOR2BX1 U297 ( .AN(a[12]), .B(n85), .Y(n179) );
  XNOR3X2 U298 ( .A(n398), .B(n358), .C(n195), .Y(c[0]) );
  XOR2X1 U299 ( .A(n286), .B(n278), .Y(n300) );
  NAND2X1 U300 ( .A(n85), .B(n97), .Y(n286) );
  OAI2BB1X1 U301 ( .A0N(n32), .A1N(n298), .B0(n297), .Y(n299) );
  XOR2X1 U302 ( .A(n153), .B(n152), .Y(n165) );
  NAND2X1 U303 ( .A(n87), .B(a[8]), .Y(n153) );
  NAND2X1 U304 ( .A(n86), .B(n16), .Y(n152) );
  XOR2X1 U305 ( .A(n146), .B(n145), .Y(n148) );
  XOR2X1 U306 ( .A(n396), .B(n397), .Y(n134) );
  XOR3X2 U307 ( .A(n422), .B(n423), .C(n384), .Y(n431) );
  XOR2X1 U308 ( .A(n421), .B(n420), .Y(n423) );
  XOR2X1 U309 ( .A(n419), .B(n418), .Y(n420) );
  XNOR3X2 U310 ( .A(n484), .B(n266), .C(n265), .Y(n302) );
  XOR3X2 U311 ( .A(n485), .B(n486), .C(n483), .Y(n266) );
  XNOR3X2 U312 ( .A(n58), .B(n451), .C(n170), .Y(n203) );
  NOR2X1 U313 ( .A(n386), .B(n388), .Y(n451) );
  XNOR2X1 U314 ( .A(n454), .B(n455), .Y(n170) );
  XOR2X1 U315 ( .A(n417), .B(n416), .Y(n418) );
  NAND2X1 U316 ( .A(n100), .B(b[9]), .Y(n443) );
  XNOR3X2 U317 ( .A(n408), .B(n361), .C(n360), .Y(n373) );
  XNOR2X1 U318 ( .A(n407), .B(n410), .Y(n360) );
  OAI2BB1X1 U319 ( .A0N(n83), .A1N(n163), .B0(n162), .Y(n164) );
  OAI21XL U320 ( .A0(n155), .A1(n176), .B0(n84), .Y(n162) );
  INVX1 U321 ( .A(n84), .Y(n154) );
  NAND2BX1 U322 ( .AN(n57), .B(n36), .Y(n381) );
  XNOR3X2 U323 ( .A(n74), .B(n77), .C(n395), .Y(n127) );
  XOR3X2 U324 ( .A(n132), .B(n131), .C(n130), .Y(n133) );
  XOR2X1 U325 ( .A(n442), .B(n441), .Y(n446) );
  NOR2X1 U326 ( .A(n386), .B(n489), .Y(n441) );
  AOI22X1 U327 ( .A0(n26), .A1(n440), .B0(n24), .B1(n439), .Y(n442) );
  OAI21XL U328 ( .A0(n24), .A1(n495), .B0(n8), .Y(n440) );
  OAI2BB1X1 U329 ( .A0N(n29), .A1N(n249), .B0(n248), .Y(n250) );
  AOI21X1 U330 ( .A0(n86), .A1(n216), .B0(n215), .Y(n217) );
  XOR3X2 U331 ( .A(n175), .B(n174), .C(n173), .Y(n182) );
  XOR2X1 U332 ( .A(n383), .B(n415), .Y(n419) );
  NAND3BX1 U333 ( .AN(n382), .B(n381), .C(n380), .Y(n383) );
  XOR2X1 U334 ( .A(n389), .B(n414), .Y(n421) );
  XOR2X1 U335 ( .A(n413), .B(n412), .Y(n414) );
  XOR3X2 U336 ( .A(n411), .B(n375), .C(n374), .Y(n389) );
  XOR2X1 U337 ( .A(n479), .B(n478), .Y(n480) );
  XOR2X1 U338 ( .A(n477), .B(n476), .Y(n478) );
  XOR2X1 U339 ( .A(n475), .B(n474), .Y(n479) );
  INVX1 U340 ( .A(n178), .Y(n181) );
  OAI21XL U341 ( .A0(n177), .A1(n176), .B0(n85), .Y(n178) );
  NOR2BX1 U342 ( .AN(n36), .B(n32), .Y(n296) );
  NOR2BX1 U343 ( .AN(a[12]), .B(n83), .Y(n139) );
  NOR2BX1 U344 ( .AN(n36), .B(n29), .Y(n247) );
  NOR2BX1 U345 ( .AN(n36), .B(n82), .Y(n111) );
  XNOR3X2 U346 ( .A(n346), .B(n343), .C(n339), .Y(n347) );
  XOR3X2 U347 ( .A(n338), .B(n337), .C(n336), .Y(n339) );
  XOR2X1 U348 ( .A(n384), .B(n500), .Y(n346) );
  XOR2X1 U349 ( .A(n459), .B(n210), .Y(n221) );
  XOR3X2 U350 ( .A(n205), .B(n204), .C(n458), .Y(n210) );
  AOI22XL U351 ( .A0(n23), .A1(n457), .B0(a[4]), .B1(n456), .Y(n459) );
  NOR2X1 U352 ( .A(n489), .B(n494), .Y(n458) );
  NAND2BXL U353 ( .AN(n87), .B(n36), .Y(n225) );
  AND2X2 U354 ( .A(n13), .B(a[3]), .Y(n151) );
  XNOR3X2 U355 ( .A(n78), .B(n79), .C(n435), .Y(n142) );
  AND2X2 U356 ( .A(n34), .B(n85), .Y(n166) );
  NAND2BXL U357 ( .AN(b[9]), .B(n37), .Y(n316) );
  XNOR2X1 U358 ( .A(n437), .B(n434), .Y(n147) );
  XNOR2X1 U359 ( .A(n449), .B(n450), .Y(n192) );
  XNOR2X1 U360 ( .A(n329), .B(n327), .Y(n330) );
  XOR2X1 U361 ( .A(n493), .B(n490), .Y(n327) );
  XNOR3X2 U362 ( .A(n326), .B(n492), .C(n361), .Y(n329) );
  INVX1 U363 ( .A(n92), .Y(n319) );
  OAI21XL U364 ( .A0(n98), .A1(n376), .B0(n8), .Y(n457) );
  OAI21XL U365 ( .A0(n21), .A1(n376), .B0(n8), .Y(n482) );
  XOR2X1 U366 ( .A(n304), .B(n303), .Y(n332) );
  NOR2BX1 U367 ( .AN(n17), .B(n489), .Y(n407) );
  NOR2X1 U368 ( .A(n386), .B(n10), .Y(n398) );
  XNOR3X2 U369 ( .A(n364), .B(n363), .C(n362), .Y(n372) );
  NAND2X1 U370 ( .A(n32), .B(a[1]), .Y(n351) );
  NAND2X1 U371 ( .A(n96), .B(n7), .Y(n352) );
  XOR2X1 U372 ( .A(n354), .B(n353), .Y(n355) );
  XOR2X1 U373 ( .A(n427), .B(n426), .Y(n428) );
  XOR2X1 U374 ( .A(n469), .B(n468), .Y(n470) );
  INVX1 U375 ( .A(n96), .Y(n386) );
  XOR2X1 U376 ( .A(n425), .B(n424), .Y(n429) );
  AOI22X1 U377 ( .A0(a[0]), .A1(n433), .B0(n26), .B1(n432), .Y(n438) );
  OAI21XL U378 ( .A0(n26), .A1(n495), .B0(n8), .Y(n433) );
  OAI21XL U379 ( .A0(n96), .A1(n10), .B0(n9), .Y(n432) );
  XOR2X1 U380 ( .A(n366), .B(n365), .Y(n367) );
  INVX1 U381 ( .A(n97), .Y(n494) );
  INVX1 U382 ( .A(b[0]), .Y(n496) );
  OAI2BB1X1 U383 ( .A0N(n82), .A1N(n126), .B0(n122), .Y(n128) );
  BUFX3 U384 ( .A(a[4]), .Y(n98) );
  BUFX3 U385 ( .A(a[6]), .Y(n100) );
  BUFX3 U386 ( .A(a[2]), .Y(n97) );
  BUFX3 U387 ( .A(a[5]), .Y(n99) );
  BUFX3 U388 ( .A(b[10]), .Y(n92) );
  BUFX3 U389 ( .A(b[11]), .Y(n95) );
  BUFX3 U390 ( .A(b[3]), .Y(n83) );
  BUFX3 U391 ( .A(b[4]), .Y(n84) );
  BUFX3 U392 ( .A(b[5]), .Y(n85) );
  BUFX3 U393 ( .A(b[6]), .Y(n86) );
  BUFX3 U394 ( .A(b[7]), .Y(n87) );
  BUFX3 U395 ( .A(b[2]), .Y(n82) );
  BUFX3 U396 ( .A(a[0]), .Y(n96) );
  OAI21XL U397 ( .A0(n107), .A1(n378), .B0(n27), .Y(n108) );
  OAI21XL U398 ( .A0(n296), .A1(n378), .B0(n29), .Y(n297) );
  OAI21XL U399 ( .A0(n179), .A1(n378), .B0(n84), .Y(n180) );
  AOI21XL U400 ( .A0(n315), .A1(n214), .B0(n213), .Y(n215) );
  OAI21XL U401 ( .A0(n111), .A1(n378), .B0(b[1]), .Y(n122) );
  AOI21XL U402 ( .A0(n315), .A1(n225), .B0(n224), .Y(n228) );
  NAND2XL U403 ( .A(n315), .B(n314), .Y(n317) );
  OAI21XL U404 ( .A0(n247), .A1(n378), .B0(n87), .Y(n248) );
  OAI21XL U405 ( .A0(n139), .A1(n378), .B0(n82), .Y(n140) );
  OAI2BB1XL U406 ( .A0N(a[12]), .A1N(n154), .B0(n315), .Y(n163) );
endmodule


module multiplier_6 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n36, n37, n38, n39, n47, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n61, n63, n64, n77, n81, n83, n84, n85,
         n86, n87, n92, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n122, n127, n128, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n202, n203, n204, n205, n210,
         n211, n212, n213, n214, n215, n216, n217, n219, n220, n221, n222,
         n239, n240, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n259, n260, n261, n262, n263, n264, n265, n266, n286, n288, n289,
         n290, n291, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n311, n314, n315, n316, n317, n318, n319, n320, n321,
         n323, n324, n325, n326, n327, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540;

  NOR2BXL U1 ( .AN(n31), .B(b[9]), .Y(n302) );
  NAND2XL U2 ( .A(b[9]), .B(n26), .Y(n265) );
  INVX1 U3 ( .A(n86), .Y(n317) );
  INVX1 U4 ( .A(n317), .Y(n2) );
  XOR2X1 U5 ( .A(n213), .B(n378), .Y(n290) );
  INVX1 U6 ( .A(n138), .Y(n334) );
  AND2X1 U7 ( .A(n14), .B(n32), .Y(n319) );
  AND2X2 U8 ( .A(n86), .B(n27), .Y(n247) );
  OAI21XL U9 ( .A0(n367), .A1(n81), .B0(n369), .Y(n141) );
  XOR3X2 U10 ( .A(n464), .B(n463), .C(n466), .Y(n494) );
  NOR2X1 U11 ( .A(n521), .B(n25), .Y(n414) );
  XNOR2X1 U12 ( .A(n138), .B(n216), .Y(n366) );
  XNOR3X2 U13 ( .A(n380), .B(n467), .C(n180), .Y(c[2]) );
  NAND2BX1 U14 ( .AN(n166), .B(n169), .Y(n170) );
  OAI2BB1X1 U15 ( .A0N(n304), .A1N(n15), .B0(n303), .Y(n305) );
  AND2X1 U16 ( .A(n81), .B(n96), .Y(n480) );
  XNOR2X1 U17 ( .A(n214), .B(n446), .Y(c[1]) );
  OAI221XL U18 ( .A0(n367), .A1(n5), .B0(n1), .B1(n7), .C0(n370), .Y(n371) );
  INVX1 U19 ( .A(n31), .Y(n1) );
  NAND3XL U20 ( .A(n163), .B(n166), .C(n168), .Y(n173) );
  XOR2X1 U21 ( .A(n493), .B(n492), .Y(c[5]) );
  XOR3X2 U22 ( .A(n354), .B(n338), .C(n353), .Y(c[10]) );
  CLKINVX3 U23 ( .A(n316), .Y(n376) );
  AOI21X1 U24 ( .A0(n316), .A1(n102), .B0(n317), .Y(n103) );
  XOR2X2 U25 ( .A(n105), .B(n58), .Y(n138) );
  AOI21X2 U26 ( .A0(n34), .A1(n104), .B0(n103), .Y(n105) );
  NOR2X1 U27 ( .A(n372), .B(n395), .Y(n373) );
  BUFX3 U28 ( .A(b[10]), .Y(n86) );
  AOI2BB2XL U29 ( .B0(b[0]), .B1(n376), .A0N(n77), .A1N(n368), .Y(n370) );
  BUFX2 U30 ( .A(n369), .Y(n77) );
  OAI21X1 U31 ( .A0(n377), .A1(n376), .B0(n375), .Y(n451) );
  NOR2X1 U32 ( .A(n262), .B(n261), .Y(n286) );
  INVX1 U33 ( .A(n213), .Y(n219) );
  INVX1 U34 ( .A(n4), .Y(n6) );
  CLKBUFXL U35 ( .A(a[12]), .Y(n31) );
  INVXL U36 ( .A(b[3]), .Y(n395) );
  INVX2 U37 ( .A(n494), .Y(n384) );
  INVX1 U38 ( .A(b[0]), .Y(n3) );
  AND2X2 U39 ( .A(b[1]), .B(n533), .Y(n4) );
  INVX1 U40 ( .A(n4), .Y(n5) );
  NAND2X1 U41 ( .A(b[0]), .B(n532), .Y(n7) );
  NAND2X1 U42 ( .A(b[0]), .B(n532), .Y(n53) );
  INVX1 U43 ( .A(n394), .Y(n8) );
  BUFX3 U44 ( .A(b[7]), .Y(n85) );
  INVX1 U45 ( .A(n190), .Y(n9) );
  INVX1 U46 ( .A(n389), .Y(n10) );
  INVX1 U47 ( .A(b[8]), .Y(n11) );
  INVX1 U48 ( .A(n11), .Y(n12) );
  INVX1 U49 ( .A(n11), .Y(n13) );
  INVX1 U50 ( .A(b[9]), .Y(n14) );
  INVX1 U51 ( .A(n14), .Y(n15) );
  INVX1 U52 ( .A(n254), .Y(n16) );
  INVX1 U53 ( .A(b[4]), .Y(n17) );
  INVXL U54 ( .A(n17), .Y(n18) );
  INVX1 U55 ( .A(n465), .Y(n19) );
  INVX1 U56 ( .A(n500), .Y(n20) );
  INVX1 U57 ( .A(a[7]), .Y(n21) );
  INVXL U58 ( .A(n21), .Y(n22) );
  INVX1 U59 ( .A(a[8]), .Y(n23) );
  INVX1 U60 ( .A(n23), .Y(n24) );
  INVX1 U61 ( .A(a[9]), .Y(n25) );
  INVX1 U62 ( .A(n25), .Y(n26) );
  INVX1 U63 ( .A(n25), .Y(n27) );
  INVX1 U64 ( .A(a[10]), .Y(n28) );
  INVX1 U65 ( .A(n28), .Y(n29) );
  INVXL U66 ( .A(n28), .Y(n30) );
  INVX1 U67 ( .A(n367), .Y(n32) );
  BUFX3 U68 ( .A(a[11]), .Y(n101) );
  OAI21XL U69 ( .A0(n100), .A1(n368), .B0(n6), .Y(n499) );
  NAND2BX4 U70 ( .AN(n101), .B(a[12]), .Y(n316) );
  INVXL U71 ( .A(n395), .Y(n33) );
  BUFX3 U72 ( .A(b[11]), .Y(n34) );
  OAI2BB1X1 U73 ( .A0N(n101), .A1N(n317), .B0(n369), .Y(n104) );
  AOI22XL U74 ( .A0(n10), .A1(n107), .B0(n34), .B1(n106), .Y(n381) );
  XNOR3X2 U75 ( .A(n47), .B(n411), .C(n323), .Y(n540) );
  NAND2XL U76 ( .A(n169), .B(n167), .Y(n174) );
  XNOR2X1 U77 ( .A(n381), .B(n360), .Y(n54) );
  INVX1 U78 ( .A(n83), .Y(n190) );
  AOI21X1 U79 ( .A0(n84), .A1(n193), .B0(n192), .Y(n212) );
  NAND2XL U80 ( .A(n97), .B(n33), .Y(n504) );
  NAND2X1 U81 ( .A(n12), .B(a[8]), .Y(n152) );
  NAND2XL U82 ( .A(n98), .B(n33), .Y(n513) );
  AOI22X1 U83 ( .A0(n22), .A1(n519), .B0(n24), .B1(n518), .Y(n523) );
  NAND2XL U84 ( .A(a[8]), .B(n83), .Y(n59) );
  NAND2XL U85 ( .A(n33), .B(a[6]), .Y(n539) );
  AND2X1 U86 ( .A(n24), .B(n81), .Y(n405) );
  INVXL U87 ( .A(n366), .Y(n179) );
  XOR3X2 U88 ( .A(n37), .B(n286), .C(n266), .Y(n36) );
  XNOR2X1 U89 ( .A(n253), .B(n252), .Y(n37) );
  NOR2XL U90 ( .A(n386), .B(n394), .Y(n418) );
  NOR2XL U91 ( .A(n388), .B(n395), .Y(n472) );
  NOR2XL U92 ( .A(n387), .B(n394), .Y(n514) );
  XOR3X2 U93 ( .A(n38), .B(n405), .C(n39), .Y(n353) );
  XOR3X2 U94 ( .A(n406), .B(n346), .C(n339), .Y(n38) );
  XNOR3X2 U95 ( .A(n352), .B(n351), .C(n350), .Y(n39) );
  NAND2XL U96 ( .A(n85), .B(n100), .Y(n398) );
  NAND2XL U97 ( .A(n98), .B(n86), .Y(n444) );
  NAND2XL U98 ( .A(n15), .B(n29), .Y(n246) );
  NAND2XL U99 ( .A(n8), .B(n97), .Y(n346) );
  NAND2XL U100 ( .A(n85), .B(n24), .Y(n453) );
  AOI22XL U101 ( .A0(n24), .A1(n535), .B0(n27), .B1(n534), .Y(n537) );
  NAND2XL U102 ( .A(n98), .B(b[9]), .Y(n400) );
  NAND2XL U103 ( .A(n99), .B(n12), .Y(n401) );
  OAI21XL U104 ( .A0(n319), .A1(n318), .B0(n86), .Y(n320) );
  INVXL U105 ( .A(n77), .Y(n318) );
  INVXL U106 ( .A(n85), .Y(n394) );
  NAND2XL U107 ( .A(n22), .B(n10), .Y(n249) );
  NAND2XL U108 ( .A(n31), .B(n10), .Y(n216) );
  NAND2BXL U109 ( .AN(b[11]), .B(a[12]), .Y(n102) );
  NAND2XL U110 ( .A(n24), .B(n86), .Y(n263) );
  NAND2XL U111 ( .A(n27), .B(n87), .Y(n47) );
  NAND2XL U112 ( .A(a[7]), .B(n15), .Y(n469) );
  OAI2BB1X1 U113 ( .A0N(n33), .A1N(n141), .B0(n140), .Y(n143) );
  NAND2XL U114 ( .A(n18), .B(n22), .Y(n416) );
  NAND2XL U115 ( .A(n97), .B(n18), .Y(n512) );
  NAND2XL U116 ( .A(n18), .B(n99), .Y(n538) );
  NAND2XL U117 ( .A(n92), .B(n15), .Y(n332) );
  NAND2XL U118 ( .A(n85), .B(n96), .Y(n331) );
  NAND2XL U119 ( .A(n30), .B(b[3]), .Y(n135) );
  NAND2XL U120 ( .A(n81), .B(n30), .Y(n422) );
  NAND2XL U121 ( .A(n100), .B(n86), .Y(n468) );
  NAND2XL U122 ( .A(n19), .B(n13), .Y(n410) );
  NAND2XL U123 ( .A(n84), .B(a[6]), .Y(n419) );
  NAND2XL U124 ( .A(n97), .B(n83), .Y(n516) );
  NAND2XL U125 ( .A(n16), .B(n96), .Y(n515) );
  NAND2XL U126 ( .A(n18), .B(n24), .Y(n423) );
  NAND2XL U127 ( .A(n98), .B(n18), .Y(n524) );
  NAND2XL U128 ( .A(n100), .B(b[9]), .Y(n457) );
  NAND2XL U129 ( .A(n13), .B(n95), .Y(n324) );
  NAND2XL U130 ( .A(n100), .B(n34), .Y(n482) );
  NAND2XL U131 ( .A(n92), .B(n8), .Y(n296) );
  NAND2XL U132 ( .A(n16), .B(n92), .Y(n495) );
  NAND2XL U133 ( .A(n98), .B(n34), .Y(n459) );
  NAND2XL U134 ( .A(n24), .B(n34), .Y(n248) );
  XOR2X1 U135 ( .A(n205), .B(n204), .Y(n210) );
  NAND2XL U136 ( .A(n83), .B(n30), .Y(n452) );
  NAND2XL U137 ( .A(a[8]), .B(n87), .Y(n300) );
  NAND2XL U138 ( .A(n26), .B(b[11]), .Y(n299) );
  NAND2XL U139 ( .A(n87), .B(n96), .Y(n146) );
  NAND2XL U140 ( .A(n97), .B(n34), .Y(n145) );
  NAND2XL U141 ( .A(a[2]), .B(n15), .Y(n409) );
  NAND2XL U142 ( .A(n29), .B(n87), .Y(n58) );
  NAND2XL U143 ( .A(n83), .B(n95), .Y(n496) );
  NAND2XL U144 ( .A(a[7]), .B(n86), .Y(n483) );
  NAND2XL U145 ( .A(n99), .B(n86), .Y(n460) );
  NAND2XL U146 ( .A(n77), .B(n220), .Y(n239) );
  NAND2BXL U147 ( .AN(n85), .B(n32), .Y(n220) );
  NAND2XL U148 ( .A(n98), .B(n16), .Y(n347) );
  NAND2XL U149 ( .A(n92), .B(n2), .Y(n348) );
  NAND2XL U150 ( .A(n15), .B(n95), .Y(n349) );
  NAND2XL U151 ( .A(n84), .B(a[7]), .Y(n399) );
  NAND2XL U152 ( .A(n85), .B(n22), .Y(n443) );
  NAND2XL U153 ( .A(n33), .B(n22), .Y(n408) );
  NAND2XL U154 ( .A(n18), .B(n100), .Y(n407) );
  NAND2XL U155 ( .A(a[5]), .B(n9), .Y(n339) );
  NAND2XL U156 ( .A(n84), .B(n29), .Y(n151) );
  OAI2BB1XL U157 ( .A0N(n101), .A1N(n190), .B0(n77), .Y(n193) );
  NAND2XL U158 ( .A(n33), .B(n27), .Y(n424) );
  NAND2XL U159 ( .A(a[7]), .B(n13), .Y(n458) );
  NAND2XL U160 ( .A(n96), .B(n18), .Y(n503) );
  NAND2XL U161 ( .A(n85), .B(n29), .Y(n195) );
  NAND2XL U162 ( .A(n12), .B(n26), .Y(n194) );
  NAND2XL U163 ( .A(n84), .B(n97), .Y(n325) );
  XNOR3X2 U164 ( .A(n381), .B(n49), .C(n380), .Y(n382) );
  NAND2XL U165 ( .A(n9), .B(n92), .Y(n49) );
  XOR3X2 U166 ( .A(n50), .B(n311), .C(n338), .Y(n314) );
  NAND2XL U167 ( .A(n16), .B(n95), .Y(n50) );
  NAND2BXL U168 ( .AN(n85), .B(n31), .Y(n259) );
  AOI22XL U169 ( .A0(a[6]), .A1(n509), .B0(n22), .B1(n508), .Y(n511) );
  XNOR3X2 U170 ( .A(n335), .B(n334), .C(n537), .Y(n336) );
  NAND2XL U171 ( .A(n87), .B(n95), .Y(n108) );
  NAND2XL U172 ( .A(b[11]), .B(n96), .Y(n109) );
  NAND2XL U173 ( .A(n86), .B(n97), .Y(n110) );
  NAND2XL U174 ( .A(n84), .B(a[8]), .Y(n63) );
  NAND2XL U175 ( .A(n27), .B(n83), .Y(n64) );
  NAND2XL U176 ( .A(n26), .B(b[4]), .Y(n61) );
  INVXL U177 ( .A(n100), .Y(n520) );
  NAND2XL U178 ( .A(n83), .B(n22), .Y(n420) );
  XNOR2XL U179 ( .A(n429), .B(n540), .Y(n430) );
  NAND2XL U180 ( .A(n92), .B(n10), .Y(n429) );
  NAND2XL U181 ( .A(n34), .B(n30), .Y(n411) );
  NAND2XL U182 ( .A(n98), .B(n87), .Y(n470) );
  NAND2XL U183 ( .A(n99), .B(b[11]), .Y(n471) );
  NAND2XL U184 ( .A(n99), .B(n15), .Y(n445) );
  NAND2XL U185 ( .A(n100), .B(n13), .Y(n442) );
  INVXL U186 ( .A(n84), .Y(n254) );
  INVXL U187 ( .A(n87), .Y(n389) );
  NAND2BXL U188 ( .AN(a[12]), .B(n101), .Y(n369) );
  AND2X1 U189 ( .A(n30), .B(b[4]), .Y(n144) );
  AND2X1 U190 ( .A(n92), .B(n18), .Y(n188) );
  AND2X1 U191 ( .A(n98), .B(n83), .Y(n326) );
  NAND2XL U192 ( .A(n77), .B(n301), .Y(n304) );
  XOR3X2 U193 ( .A(n52), .B(n306), .C(n305), .Y(n51) );
  NAND2XL U194 ( .A(n30), .B(n86), .Y(n52) );
  AND2X1 U195 ( .A(n22), .B(n81), .Y(n536) );
  INVXL U196 ( .A(n101), .Y(n367) );
  XOR2X1 U197 ( .A(n456), .B(n455), .Y(n464) );
  XOR2X1 U198 ( .A(n454), .B(n453), .Y(n455) );
  NAND2XL U199 ( .A(n84), .B(n27), .Y(n454) );
  NAND2XL U200 ( .A(n99), .B(n87), .Y(n203) );
  NAND2XL U201 ( .A(b[9]), .B(a[8]), .Y(n202) );
  NAND2XL U202 ( .A(n13), .B(n96), .Y(n351) );
  NAND2XL U203 ( .A(n92), .B(n34), .Y(n362) );
  NAND2XL U204 ( .A(n95), .B(b[10]), .Y(n361) );
  NAND2XL U205 ( .A(a[6]), .B(n9), .Y(n357) );
  NAND2XL U206 ( .A(a[5]), .B(n16), .Y(n358) );
  NAND2XL U207 ( .A(n20), .B(n8), .Y(n359) );
  NAND2XL U208 ( .A(n19), .B(n15), .Y(n432) );
  NAND2XL U209 ( .A(n18), .B(a[1]), .Y(n488) );
  NAND2XL U210 ( .A(a[1]), .B(n34), .Y(n434) );
  AND2X1 U211 ( .A(n13), .B(a[0]), .Y(n530) );
  NAND2XL U212 ( .A(a[2]), .B(b[10]), .Y(n435) );
  NAND2XL U213 ( .A(n20), .B(n13), .Y(n433) );
  NAND2XL U214 ( .A(n77), .B(n127), .Y(n132) );
  NAND2BXL U215 ( .AN(b[1]), .B(n101), .Y(n127) );
  INVXL U216 ( .A(b[1]), .Y(n368) );
  XOR2X1 U217 ( .A(n57), .B(n384), .Y(n288) );
  XOR2X1 U218 ( .A(n138), .B(n381), .Y(n354) );
  XOR2X1 U219 ( .A(n540), .B(n51), .Y(n356) );
  XNOR3X2 U220 ( .A(n179), .B(n178), .C(n380), .Y(n214) );
  XOR3X2 U221 ( .A(n265), .B(n264), .C(n263), .Y(n266) );
  XOR3X2 U222 ( .A(n356), .B(n530), .C(n531), .Y(c[8]) );
  XNOR3X2 U223 ( .A(n179), .B(n219), .C(n178), .Y(n181) );
  XOR2X1 U224 ( .A(n298), .B(n51), .Y(n338) );
  XNOR2X1 U225 ( .A(n494), .B(n381), .Y(n180) );
  XOR3X2 U226 ( .A(n514), .B(n36), .C(n385), .Y(n396) );
  XNOR3X2 U227 ( .A(n219), .B(n507), .C(n217), .Y(n289) );
  XOR2X1 U228 ( .A(n216), .B(n497), .Y(n217) );
  XOR2X1 U229 ( .A(n506), .B(n505), .Y(n507) );
  XOR2X1 U230 ( .A(n496), .B(n495), .Y(n497) );
  XNOR3X2 U231 ( .A(n215), .B(n290), .C(n214), .Y(c[4]) );
  XNOR3X2 U232 ( .A(n54), .B(n55), .C(n56), .Y(n363) );
  XNOR2X1 U233 ( .A(n409), .B(n410), .Y(n55) );
  XOR3X2 U234 ( .A(n416), .B(n362), .C(n361), .Y(n56) );
  INVX1 U235 ( .A(n216), .Y(n360) );
  INVX1 U236 ( .A(n385), .Y(n378) );
  XOR2X1 U237 ( .A(n289), .B(n288), .Y(c[6]) );
  XOR2X1 U238 ( .A(n439), .B(n438), .Y(c[12]) );
  XNOR2X1 U239 ( .A(n298), .B(n36), .Y(n57) );
  XOR2X1 U240 ( .A(n529), .B(n528), .Y(n531) );
  XOR2X1 U241 ( .A(n527), .B(n526), .Y(n528) );
  XOR2X1 U242 ( .A(n396), .B(n517), .Y(n529) );
  XOR2X1 U243 ( .A(n525), .B(n524), .Y(n526) );
  INVX1 U244 ( .A(n168), .Y(n169) );
  XOR2X1 U245 ( .A(n477), .B(n472), .Y(n182) );
  XOR2X1 U246 ( .A(n476), .B(n475), .Y(n477) );
  NOR2X1 U247 ( .A(n387), .B(n521), .Y(n475) );
  XOR2X1 U248 ( .A(n315), .B(n314), .Y(c[7]) );
  XNOR3X2 U249 ( .A(n182), .B(n181), .C(n180), .Y(c[3]) );
  XNOR3X2 U250 ( .A(n337), .B(n57), .C(n336), .Y(c[9]) );
  XNOR3X2 U251 ( .A(n365), .B(n364), .C(n363), .Y(c[11]) );
  NOR2X1 U252 ( .A(n521), .B(n386), .Y(n510) );
  OAI21XL U253 ( .A0(n34), .A1(n367), .B0(n77), .Y(n107) );
  NAND2BXL U254 ( .AN(n84), .B(a[12]), .Y(n191) );
  OAI21XL U255 ( .A0(n27), .A1(n532), .B0(n6), .Y(n535) );
  OAI21XL U256 ( .A0(n24), .A1(n3), .B0(n53), .Y(n534) );
  OAI2BB1X1 U257 ( .A0N(n101), .A1N(b[4]), .B0(n395), .Y(n375) );
  MXI2X1 U258 ( .A(n374), .B(n373), .S0(b[4]), .Y(n377) );
  INVXL U259 ( .A(a[12]), .Y(n374) );
  AOI22X1 U260 ( .A0(n96), .A1(n474), .B0(n97), .B1(n473), .Y(n476) );
  OAI21XL U261 ( .A0(n97), .A1(n368), .B0(n6), .Y(n474) );
  OAI21XL U262 ( .A0(n96), .A1(n3), .B0(n7), .Y(n473) );
  AOI22X1 U263 ( .A0(n30), .A1(n404), .B0(n27), .B1(n403), .Y(n406) );
  OAI21XL U264 ( .A0(n30), .A1(n368), .B0(n5), .Y(n403) );
  OAI21XL U265 ( .A0(n27), .A1(n3), .B0(n53), .Y(n404) );
  OAI21XL U266 ( .A0(n165), .A1(n372), .B0(n83), .Y(n166) );
  NOR2BX1 U267 ( .AN(n101), .B(b[4]), .Y(n165) );
  AOI21X1 U268 ( .A0(n77), .A1(n260), .B0(n394), .Y(n261) );
  NAND2BX1 U269 ( .AN(n84), .B(n101), .Y(n260) );
  OAI2BB1X1 U270 ( .A0N(n15), .A1N(n321), .B0(n320), .Y(n323) );
  OAI21XL U271 ( .A0(n24), .A1(n368), .B0(n6), .Y(n519) );
  OAI21XL U272 ( .A0(n20), .A1(n368), .B0(n6), .Y(n479) );
  OAI21XL U273 ( .A0(n22), .A1(n368), .B0(n6), .Y(n509) );
  OAI21XL U274 ( .A0(n32), .A1(n368), .B0(n6), .Y(n413) );
  OAI21XL U275 ( .A0(n99), .A1(n3), .B0(n53), .Y(n498) );
  OAI21XL U276 ( .A0(n22), .A1(n3), .B0(n7), .Y(n518) );
  OAI21XL U277 ( .A0(n95), .A1(n3), .B0(n7), .Y(n447) );
  OAI21XL U278 ( .A0(n19), .A1(n533), .B0(n53), .Y(n478) );
  AOI22X1 U279 ( .A0(n20), .A1(n485), .B0(a[5]), .B1(n484), .Y(n486) );
  OAI21XL U280 ( .A0(a[5]), .A1(n368), .B0(n6), .Y(n485) );
  OAI21XL U281 ( .A0(n98), .A1(n533), .B0(n7), .Y(n484) );
  OAI21XL U282 ( .A0(a[6]), .A1(n3), .B0(n53), .Y(n508) );
  OAI21XL U283 ( .A0(n30), .A1(n3), .B0(n53), .Y(n412) );
  INVX1 U284 ( .A(n81), .Y(n521) );
  XOR2X1 U285 ( .A(n150), .B(n149), .Y(n380) );
  XNOR3X2 U286 ( .A(n444), .B(n148), .C(n147), .Y(n149) );
  XNOR3X2 U287 ( .A(n144), .B(n143), .C(n142), .Y(n150) );
  OAI21XL U288 ( .A0(n302), .A1(n376), .B0(n13), .Y(n303) );
  XNOR3X2 U289 ( .A(n212), .B(n211), .C(n210), .Y(n385) );
  XNOR2X1 U290 ( .A(n483), .B(n482), .Y(n211) );
  XOR2X1 U291 ( .A(n137), .B(n136), .Y(n178) );
  XNOR3X2 U292 ( .A(n398), .B(n122), .C(n111), .Y(n137) );
  XNOR3X2 U293 ( .A(n135), .B(n134), .C(n133), .Y(n136) );
  XOR3X2 U294 ( .A(n153), .B(n152), .C(n151), .Y(n168) );
  NAND2X1 U295 ( .A(n85), .B(n26), .Y(n153) );
  XOR2X1 U296 ( .A(n177), .B(n176), .Y(n213) );
  XNOR3X2 U297 ( .A(n468), .B(n469), .C(n175), .Y(n176) );
  NAND3X1 U298 ( .A(n174), .B(n173), .C(n170), .Y(n177) );
  XOR2X1 U299 ( .A(n251), .B(n250), .Y(n298) );
  XOR2X1 U300 ( .A(n249), .B(n248), .Y(n250) );
  XNOR3X2 U301 ( .A(n247), .B(n246), .C(n240), .Y(n251) );
  NOR2X1 U302 ( .A(n389), .B(n465), .Y(n466) );
  INVX1 U303 ( .A(n97), .Y(n465) );
  NAND2X1 U304 ( .A(n100), .B(n87), .Y(n264) );
  NOR2BX1 U305 ( .AN(n31), .B(n13), .Y(n221) );
  NOR2BX1 U306 ( .AN(n31), .B(b[3]), .Y(n139) );
  NOR2BX1 U307 ( .AN(a[12]), .B(n81), .Y(n128) );
  OAI21XL U308 ( .A0(n139), .A1(n376), .B0(n81), .Y(n140) );
  NAND2X1 U309 ( .A(a[7]), .B(b[11]), .Y(n252) );
  XOR2X1 U310 ( .A(n300), .B(n299), .Y(n306) );
  XNOR2X1 U311 ( .A(n195), .B(n194), .Y(n205) );
  XOR2X1 U312 ( .A(n504), .B(n503), .Y(n505) );
  XOR3X2 U313 ( .A(n384), .B(n383), .C(n382), .Y(n492) );
  XOR2X1 U314 ( .A(n378), .B(n36), .Y(n383) );
  XNOR3X2 U315 ( .A(n402), .B(n354), .C(n178), .Y(c[0]) );
  NOR2X1 U316 ( .A(n388), .B(n3), .Y(n402) );
  XOR2X1 U317 ( .A(n297), .B(n296), .Y(n311) );
  NAND2X1 U318 ( .A(n9), .B(n96), .Y(n297) );
  XOR2X1 U319 ( .A(n450), .B(n449), .Y(n467) );
  NOR2X1 U320 ( .A(n388), .B(n521), .Y(n449) );
  AOI22X1 U321 ( .A0(n95), .A1(n448), .B0(a[2]), .B1(n447), .Y(n450) );
  OAI21XL U322 ( .A0(a[2]), .A1(n368), .B0(n6), .Y(n448) );
  XOR2X1 U323 ( .A(n400), .B(n401), .Y(n122) );
  XOR2X1 U324 ( .A(n146), .B(n145), .Y(n148) );
  XNOR3X2 U325 ( .A(n511), .B(n291), .C(n290), .Y(n315) );
  XOR3X2 U326 ( .A(n512), .B(n513), .C(n510), .Y(n291) );
  XOR2X1 U327 ( .A(n203), .B(n202), .Y(n204) );
  XOR2X1 U328 ( .A(n462), .B(n461), .Y(n463) );
  XOR2X1 U329 ( .A(n458), .B(n457), .Y(n462) );
  XOR2X1 U330 ( .A(n460), .B(n459), .Y(n461) );
  XOR2X1 U331 ( .A(n426), .B(n425), .Y(n427) );
  XOR2X1 U332 ( .A(n424), .B(n423), .Y(n425) );
  XOR2X1 U333 ( .A(n371), .B(n422), .Y(n426) );
  NAND2BXL U334 ( .AN(n12), .B(n32), .Y(n301) );
  NAND2X1 U335 ( .A(n12), .B(n29), .Y(n253) );
  XNOR3X2 U336 ( .A(n415), .B(n356), .C(n355), .Y(n365) );
  XNOR2X1 U337 ( .A(n414), .B(n417), .Y(n355) );
  AOI22XL U338 ( .A0(n30), .A1(n413), .B0(n32), .B1(n412), .Y(n415) );
  NAND2X1 U339 ( .A(n33), .B(n24), .Y(n417) );
  XNOR3X2 U340 ( .A(n330), .B(n327), .C(n540), .Y(n337) );
  XOR2X1 U341 ( .A(n325), .B(n324), .Y(n330) );
  XOR2X1 U342 ( .A(n536), .B(n326), .Y(n327) );
  XNOR3X2 U343 ( .A(n59), .B(n61), .C(n399), .Y(n133) );
  XNOR3X2 U344 ( .A(n63), .B(n64), .C(n443), .Y(n142) );
  XOR3X2 U345 ( .A(n538), .B(n539), .C(n333), .Y(n335) );
  XNOR3X2 U346 ( .A(n110), .B(n109), .C(n108), .Y(n111) );
  OAI2BB1X1 U347 ( .A0N(n13), .A1N(n239), .B0(n222), .Y(n240) );
  OAI21XL U348 ( .A0(n221), .A1(n376), .B0(n85), .Y(n222) );
  XOR2X1 U349 ( .A(n502), .B(n501), .Y(n506) );
  NOR2X1 U350 ( .A(n521), .B(n500), .Y(n501) );
  AOI22X1 U351 ( .A0(n99), .A1(n499), .B0(n100), .B1(n498), .Y(n502) );
  INVX1 U352 ( .A(n98), .Y(n500) );
  XOR2X1 U353 ( .A(n523), .B(n522), .Y(n527) );
  NOR2X1 U354 ( .A(n521), .B(n520), .Y(n522) );
  XOR2X1 U355 ( .A(n452), .B(n451), .Y(n456) );
  XOR2X1 U356 ( .A(n431), .B(n430), .Y(n439) );
  XOR2X1 U357 ( .A(n428), .B(n427), .Y(n431) );
  XOR2X1 U358 ( .A(n397), .B(n421), .Y(n428) );
  XOR2X1 U359 ( .A(n420), .B(n419), .Y(n421) );
  XOR2X1 U360 ( .A(n366), .B(n418), .Y(n397) );
  XOR2X1 U361 ( .A(n491), .B(n490), .Y(n493) );
  XOR2X1 U362 ( .A(n489), .B(n488), .Y(n490) );
  XOR2X1 U363 ( .A(n487), .B(n486), .Y(n491) );
  NAND2X1 U364 ( .A(a[2]), .B(n33), .Y(n489) );
  INVX1 U365 ( .A(n163), .Y(n167) );
  OAI21XL U366 ( .A0(n162), .A1(n376), .B0(n18), .Y(n163) );
  NOR2BX1 U367 ( .AN(n31), .B(n83), .Y(n162) );
  XOR2X1 U368 ( .A(n481), .B(n189), .Y(n215) );
  XOR3X2 U369 ( .A(n188), .B(n187), .C(n480), .Y(n189) );
  AOI22X1 U370 ( .A0(n19), .A1(n479), .B0(n20), .B1(n478), .Y(n481) );
  INVX1 U371 ( .A(n164), .Y(n372) );
  NAND2BX1 U372 ( .AN(a[12]), .B(n101), .Y(n164) );
  XNOR2X1 U373 ( .A(n470), .B(n471), .Y(n175) );
  XNOR2X1 U374 ( .A(n445), .B(n442), .Y(n147) );
  AOI22X1 U375 ( .A0(a[0]), .A1(n441), .B0(a[1]), .B1(n440), .Y(n446) );
  OAI21XL U376 ( .A0(a[1]), .A1(n532), .B0(n6), .Y(n441) );
  OAI21XL U377 ( .A0(n92), .A1(n3), .B0(n7), .Y(n440) );
  XOR2X1 U378 ( .A(n516), .B(n515), .Y(n517) );
  XOR2X1 U379 ( .A(n437), .B(n436), .Y(n438) );
  XOR2X1 U380 ( .A(n433), .B(n432), .Y(n437) );
  XOR2X1 U381 ( .A(n435), .B(n434), .Y(n436) );
  AND2X2 U382 ( .A(n33), .B(n95), .Y(n187) );
  NAND2X1 U383 ( .A(n99), .B(n33), .Y(n525) );
  NAND2X1 U384 ( .A(n19), .B(n81), .Y(n487) );
  XOR3X2 U385 ( .A(n349), .B(n348), .C(n347), .Y(n350) );
  XNOR3X2 U386 ( .A(n359), .B(n358), .C(n357), .Y(n364) );
  INVX1 U387 ( .A(n92), .Y(n388) );
  XOR2X1 U388 ( .A(n332), .B(n331), .Y(n333) );
  XOR2X1 U389 ( .A(n408), .B(n407), .Y(n352) );
  INVX1 U390 ( .A(n95), .Y(n387) );
  INVX1 U391 ( .A(n99), .Y(n386) );
  OAI2BB1X1 U392 ( .A0N(n81), .A1N(n132), .B0(n131), .Y(n134) );
  OAI21XL U393 ( .A0(n128), .A1(n376), .B0(b[1]), .Y(n131) );
  BUFX3 U394 ( .A(a[3]), .Y(n97) );
  BUFX3 U395 ( .A(a[6]), .Y(n100) );
  BUFX3 U396 ( .A(a[2]), .Y(n96) );
  BUFX3 U397 ( .A(a[4]), .Y(n98) );
  BUFX3 U398 ( .A(a[5]), .Y(n99) );
  BUFX3 U399 ( .A(b[6]), .Y(n84) );
  BUFX3 U400 ( .A(a[1]), .Y(n95) );
  BUFX3 U401 ( .A(b[12]), .Y(n87) );
  BUFX3 U402 ( .A(b[5]), .Y(n83) );
  INVX1 U403 ( .A(b[0]), .Y(n533) );
  INVX1 U404 ( .A(b[1]), .Y(n532) );
  BUFX3 U405 ( .A(b[2]), .Y(n81) );
  BUFX3 U406 ( .A(a[0]), .Y(n92) );
  OAI21XL U407 ( .A0(n87), .A1(n374), .B0(n316), .Y(n106) );
  OAI2BB1X1 U408 ( .A0N(n31), .A1N(n317), .B0(n316), .Y(n321) );
  AOI21X1 U409 ( .A0(n316), .A1(n191), .B0(n190), .Y(n192) );
  AOI21X1 U410 ( .A0(n316), .A1(n259), .B0(n254), .Y(n262) );
endmodule


module multiplier_5 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n49, n50, n51, n52, n53,
         n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n74, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n92, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n119, n122, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n202,
         n203, n204, n205, n210, n211, n212, n213, n214, n215, n216, n217,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n230,
         n233, n234, n235, n236, n237, n238, n239, n240, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n259, n260, n261, n262, n263,
         n264, n265, n266, n278, n286, n288, n289, n290, n291, n292, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n343, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494;

  NAND2XL U1 ( .A(n20), .B(b[3]), .Y(n459) );
  NAND2XL U2 ( .A(b[3]), .B(a[6]), .Y(n494) );
  NAND2XL U3 ( .A(a[0]), .B(b[5]), .Y(n239) );
  NAND2XL U4 ( .A(a[4]), .B(b[5]), .Y(n333) );
  XOR2X1 U5 ( .A(n154), .B(n153), .Y(n175) );
  NOR2X1 U6 ( .A(n30), .B(n37), .Y(n296) );
  OAI21XL U7 ( .A0(n96), .A1(n32), .B0(n376), .Y(n250) );
  OAI21XL U8 ( .A0(n97), .A1(n37), .B0(n317), .Y(n318) );
  OAI21XL U9 ( .A0(n32), .A1(n29), .B0(n376), .Y(n1) );
  INVX1 U10 ( .A(n1), .Y(n52) );
  NOR2BX1 U11 ( .AN(n102), .B(n480), .Y(n465) );
  NOR2X1 U12 ( .A(n37), .B(n92), .Y(n187) );
  NOR2X1 U13 ( .A(n32), .B(n87), .Y(n181) );
  NOR2BX1 U14 ( .AN(n104), .B(n480), .Y(n481) );
  OAI21XL U15 ( .A0(n2), .A1(n322), .B0(n323), .Y(n324) );
  INVX1 U16 ( .A(n321), .Y(n2) );
  OR2X2 U17 ( .A(n188), .B(n189), .Y(n190) );
  NOR2X1 U18 ( .A(n18), .B(n480), .Y(n446) );
  AOI211X1 U19 ( .A0(n318), .A1(n30), .B0(n323), .C0(n31), .Y(n3) );
  INVX1 U20 ( .A(n3), .Y(n326) );
  NOR2X1 U21 ( .A(n16), .B(n37), .Y(n248) );
  OAI21XL U22 ( .A0(n377), .A1(n106), .B0(n97), .Y(n107) );
  OR2X2 U23 ( .A(n189), .B(n182), .Y(n192) );
  XOR3X2 U24 ( .A(n369), .B(n401), .C(n368), .Y(n370) );
  OAI221XL U25 ( .A0(n32), .A1(n9), .B0(n487), .B1(n37), .C0(n378), .Y(n380)
         );
  NAND3X1 U26 ( .A(n182), .B(n188), .C(n189), .Y(n191) );
  XNOR2X1 U27 ( .A(n221), .B(n430), .Y(c[1]) );
  CLKINVX3 U28 ( .A(n317), .Y(n377) );
  NAND2BX1 U29 ( .AN(a[11]), .B(a[12]), .Y(n317) );
  INVX1 U30 ( .A(n373), .Y(n141) );
  XOR2X1 U31 ( .A(n413), .B(n412), .Y(n415) );
  XNOR3X2 U32 ( .A(n238), .B(n237), .C(n236), .Y(n4) );
  XNOR3X2 U33 ( .A(n50), .B(n51), .C(n299), .Y(n5) );
  AND2X2 U34 ( .A(b[1]), .B(n488), .Y(n6) );
  INVX1 U35 ( .A(n487), .Y(n7) );
  INVXL U36 ( .A(n7), .Y(n8) );
  INVX1 U37 ( .A(n6), .Y(n9) );
  INVXL U38 ( .A(n6), .Y(n10) );
  INVX1 U39 ( .A(b[0]), .Y(n11) );
  INVX1 U40 ( .A(b[0]), .Y(n488) );
  BUFX3 U41 ( .A(n376), .Y(n85) );
  INVX1 U42 ( .A(n384), .Y(n12) );
  BUFX3 U43 ( .A(n99), .Y(n13) );
  INVX1 U44 ( .A(n225), .Y(n14) );
  INVX1 U45 ( .A(b[8]), .Y(n15) );
  INVX1 U46 ( .A(n15), .Y(n16) );
  INVX1 U47 ( .A(n111), .Y(n17) );
  OAI2BB1X2 U48 ( .A0N(n98), .A1N(n108), .B0(n107), .Y(n110) );
  INVX1 U49 ( .A(a[1]), .Y(n18) );
  INVX1 U50 ( .A(n18), .Y(n19) );
  INVX1 U51 ( .A(n485), .Y(n20) );
  INVX1 U52 ( .A(a[3]), .Y(n21) );
  INVXL U53 ( .A(n21), .Y(n22) );
  INVX1 U54 ( .A(a[7]), .Y(n23) );
  INVXL U55 ( .A(n23), .Y(n24) );
  INVX1 U56 ( .A(a[8]), .Y(n25) );
  INVX1 U57 ( .A(n25), .Y(n26) );
  INVX1 U58 ( .A(n399), .Y(n27) );
  INVX1 U59 ( .A(b[9]), .Y(n28) );
  INVX1 U60 ( .A(n28), .Y(n29) );
  INVXL U61 ( .A(n28), .Y(n30) );
  INVX1 U62 ( .A(n320), .Y(n31) );
  INVX1 U63 ( .A(a[11]), .Y(n32) );
  INVXL U64 ( .A(n32), .Y(n33) );
  NAND2BX1 U65 ( .AN(a[12]), .B(a[11]), .Y(n376) );
  XOR2X2 U66 ( .A(n195), .B(n194), .Y(n262) );
  XOR2X2 U67 ( .A(n202), .B(n175), .Y(n77) );
  INVX1 U68 ( .A(a[10]), .Y(n34) );
  INVX1 U69 ( .A(n34), .Y(n35) );
  INVXL U70 ( .A(n34), .Y(n36) );
  AND2X1 U71 ( .A(n35), .B(n99), .Y(n109) );
  INVX1 U72 ( .A(a[12]), .Y(n37) );
  INVXL U73 ( .A(n37), .Y(n38) );
  OAI2BB1XL U74 ( .A0N(n33), .A1N(n111), .B0(n85), .Y(n126) );
  XOR2X1 U75 ( .A(n262), .B(n67), .Y(n266) );
  AOI2BB2XL U76 ( .B0(b[0]), .B1(n377), .A0N(n85), .A1N(n375), .Y(n378) );
  XOR2XL U77 ( .A(n289), .B(n5), .Y(n359) );
  XNOR3X2 U78 ( .A(n173), .B(n39), .C(n49), .Y(n263) );
  XNOR3X2 U79 ( .A(n155), .B(n437), .C(n79), .Y(n39) );
  XNOR3X2 U80 ( .A(n170), .B(n169), .C(n168), .Y(n49) );
  XOR2X1 U81 ( .A(n77), .B(n438), .Y(c[2]) );
  NAND2XL U82 ( .A(n102), .B(n97), .Y(n428) );
  AOI22XL U83 ( .A0(n20), .A1(n445), .B0(n22), .B1(n444), .Y(n447) );
  AOI22XL U84 ( .A0(n26), .A1(n490), .B0(n27), .B1(n489), .Y(n492) );
  NAND2XL U85 ( .A(n96), .B(n104), .Y(n386) );
  AOI22XL U86 ( .A0(n36), .A1(n392), .B0(n27), .B1(n391), .Y(n393) );
  NAND2XL U87 ( .A(n85), .B(n142), .Y(n145) );
  NAND2XL U88 ( .A(n87), .B(a[6]), .Y(n394) );
  NAND2XL U89 ( .A(b[8]), .B(n36), .Y(n234) );
  NAND2XL U90 ( .A(n30), .B(n36), .Y(n252) );
  NAND2XL U91 ( .A(n103), .B(n97), .Y(n437) );
  NAND2BXL U92 ( .AN(n95), .B(n38), .Y(n215) );
  NAND2XL U93 ( .A(n105), .B(n99), .Y(n316) );
  NAND2XL U94 ( .A(n96), .B(a[8]), .Y(n163) );
  NAND2XL U95 ( .A(n95), .B(n105), .Y(n162) );
  NAND2XL U96 ( .A(n99), .B(n101), .Y(n150) );
  NAND2XL U97 ( .A(a[3]), .B(n98), .Y(n149) );
  NAND2XL U98 ( .A(n103), .B(b[8]), .Y(n389) );
  INVXL U99 ( .A(n95), .Y(n225) );
  NOR2X1 U100 ( .A(n230), .B(n228), .Y(n237) );
  AOI21XL U101 ( .A0(n85), .A1(n227), .B0(n384), .Y(n228) );
  NAND2XL U102 ( .A(n36), .B(n97), .Y(n50) );
  XNOR2X1 U103 ( .A(n291), .B(n290), .Y(n51) );
  NAND2XL U104 ( .A(n38), .B(n99), .Y(n363) );
  NAND2XL U105 ( .A(n24), .B(n13), .Y(n259) );
  NAND2XL U106 ( .A(n85), .B(n292), .Y(n298) );
  NOR2BXL U107 ( .AN(n38), .B(n13), .Y(n119) );
  NAND2XL U108 ( .A(a[7]), .B(n17), .Y(n233) );
  NOR2BXL U109 ( .AN(a[12]), .B(n98), .Y(n106) );
  NAND2XL U110 ( .A(n104), .B(n31), .Y(n439) );
  NAND2XL U111 ( .A(n29), .B(n105), .Y(n235) );
  NAND2XL U112 ( .A(n22), .B(b[4]), .Y(n476) );
  NAND2XL U113 ( .A(b[4]), .B(n19), .Y(n458) );
  INVXL U114 ( .A(n96), .Y(n384) );
  NAND2XL U115 ( .A(n103), .B(n99), .Y(n212) );
  NAND2XL U116 ( .A(n95), .B(n104), .Y(n405) );
  NAND2XL U117 ( .A(n104), .B(n16), .Y(n426) );
  NAND2XL U118 ( .A(n103), .B(n29), .Y(n429) );
  NAND2XL U119 ( .A(n86), .B(n27), .Y(n409) );
  NAND2XL U120 ( .A(n87), .B(n26), .Y(n408) );
  NAND2XL U121 ( .A(a[7]), .B(n97), .Y(n453) );
  NAND2XL U122 ( .A(n105), .B(n98), .Y(n290) );
  NAND2XL U123 ( .A(n26), .B(n17), .Y(n254) );
  NAND2XL U124 ( .A(n104), .B(n99), .Y(n223) );
  NAND2XL U125 ( .A(a[7]), .B(b[8]), .Y(n436) );
  NAND2XL U126 ( .A(n95), .B(n100), .Y(n460) );
  NAND2XL U127 ( .A(n96), .B(n36), .Y(n213) );
  NAND2XL U128 ( .A(n26), .B(n97), .Y(n224) );
  NAND2XL U129 ( .A(n104), .B(n98), .Y(n452) );
  NAND2XL U130 ( .A(n100), .B(n17), .Y(n364) );
  NAND2XL U131 ( .A(a[8]), .B(n99), .Y(n291) );
  INVXL U132 ( .A(n103), .Y(n382) );
  AOI22XL U133 ( .A0(n22), .A1(n449), .B0(n102), .B1(n448), .Y(n451) );
  XNOR3X2 U134 ( .A(n53), .B(n54), .C(n219), .Y(n220) );
  NAND2XL U135 ( .A(n29), .B(n26), .Y(n53) );
  NAND2XL U136 ( .A(n16), .B(n105), .Y(n54) );
  NAND2XL U137 ( .A(n96), .B(a[7]), .Y(n427) );
  NAND2XL U138 ( .A(n95), .B(a[7]), .Y(n387) );
  NAND2XL U139 ( .A(b[3]), .B(n26), .Y(n403) );
  INVXL U140 ( .A(n105), .Y(n399) );
  NAND2XL U141 ( .A(n95), .B(n35), .Y(n177) );
  NAND2XL U142 ( .A(n96), .B(n22), .Y(n354) );
  NAND2XL U143 ( .A(n103), .B(n92), .Y(n353) );
  NAND2XL U144 ( .A(a[3]), .B(n86), .Y(n468) );
  NAND2XL U145 ( .A(n101), .B(n87), .Y(n467) );
  NAND2BXL U146 ( .AN(n95), .B(a[11]), .Y(n227) );
  XOR3X2 U147 ( .A(n55), .B(n402), .C(n365), .Y(n366) );
  NAND2XL U148 ( .A(a[1]), .B(n31), .Y(n55) );
  XOR3X2 U149 ( .A(n57), .B(n300), .C(n359), .Y(n301) );
  NAND2XL U150 ( .A(n14), .B(n19), .Y(n57) );
  XOR2X1 U151 ( .A(n58), .B(n59), .Y(n413) );
  XNOR3X2 U152 ( .A(n404), .B(n374), .C(n373), .Y(n58) );
  XNOR2X1 U153 ( .A(n406), .B(n405), .Y(n59) );
  NAND2XL U154 ( .A(n100), .B(n13), .Y(n414) );
  XOR3X2 U155 ( .A(n60), .B(n483), .C(n368), .Y(n328) );
  NAND2XL U156 ( .A(n100), .B(n16), .Y(n60) );
  XOR3X2 U157 ( .A(n61), .B(n352), .C(n351), .Y(n356) );
  NAND2XL U158 ( .A(n26), .B(b[2]), .Y(n61) );
  XOR3X2 U159 ( .A(n62), .B(n396), .C(n84), .Y(n367) );
  NAND2XL U160 ( .A(a[3]), .B(n16), .Y(n62) );
  NAND2XL U161 ( .A(n13), .B(a[1]), .Y(n134) );
  NAND2XL U162 ( .A(n98), .B(n101), .Y(n135) );
  NAND2XL U163 ( .A(n97), .B(a[3]), .Y(n136) );
  NAND2XL U164 ( .A(n95), .B(a[8]), .Y(n82) );
  NAND2XL U165 ( .A(n105), .B(n92), .Y(n83) );
  NAND2XL U166 ( .A(a[8]), .B(n92), .Y(n80) );
  NAND2XL U167 ( .A(n105), .B(n87), .Y(n81) );
  NAND2XL U168 ( .A(n16), .B(n19), .Y(n343) );
  OAI2BB1X1 U169 ( .A0N(a[11]), .A1N(n320), .B0(n376), .Y(n108) );
  NAND2BXL U170 ( .AN(b[2]), .B(a[11]), .Y(n142) );
  NAND2BXL U171 ( .AN(b[8]), .B(n33), .Y(n292) );
  NAND2XL U172 ( .A(n102), .B(n99), .Y(n441) );
  NAND2XL U173 ( .A(n103), .B(n98), .Y(n442) );
  INVX1 U174 ( .A(n482), .Y(n306) );
  AOI22XL U175 ( .A0(n24), .A1(n479), .B0(n26), .B1(n478), .Y(n482) );
  AOI22XL U176 ( .A0(n36), .A1(n398), .B0(n33), .B1(n397), .Y(n401) );
  NOR2XL U177 ( .A(n383), .B(n11), .Y(n390) );
  AND2X1 U178 ( .A(n102), .B(n98), .Y(n79) );
  NAND2XL U179 ( .A(a[5]), .B(b[3]), .Y(n484) );
  AND2X1 U180 ( .A(n35), .B(n87), .Y(n148) );
  AND2X1 U181 ( .A(n36), .B(n86), .Y(n133) );
  AND2X1 U182 ( .A(n105), .B(n97), .Y(n253) );
  AND2X1 U183 ( .A(n14), .B(n101), .Y(n314) );
  AND2X1 U184 ( .A(n100), .B(n87), .Y(n210) );
  INVXL U185 ( .A(n98), .Y(n111) );
  NAND2XL U186 ( .A(n12), .B(n101), .Y(n337) );
  NAND2XL U187 ( .A(n103), .B(n14), .Y(n361) );
  NAND2XL U188 ( .A(n14), .B(n22), .Y(n336) );
  NAND2XL U189 ( .A(b[4]), .B(a[5]), .Y(n493) );
  NAND2XL U190 ( .A(a[4]), .B(n14), .Y(n349) );
  NAND2XL U191 ( .A(n12), .B(n19), .Y(n303) );
  NAND2XL U192 ( .A(n22), .B(b[2]), .Y(n457) );
  NAND2XL U193 ( .A(n16), .B(n101), .Y(n350) );
  NAND2XL U194 ( .A(b[5]), .B(n22), .Y(n304) );
  NAND2XL U195 ( .A(a[4]), .B(n12), .Y(n360) );
  NAND2XL U196 ( .A(n20), .B(n31), .Y(n419) );
  NAND2XL U197 ( .A(n19), .B(n17), .Y(n418) );
  NAND2XL U198 ( .A(a[4]), .B(n16), .Y(n417) );
  NAND2XL U199 ( .A(n22), .B(n30), .Y(n416) );
  NAND2XL U200 ( .A(n85), .B(n127), .Y(n130) );
  INVX1 U201 ( .A(b[1]), .Y(n486) );
  NAND2XL U202 ( .A(b[0]), .B(n486), .Y(n487) );
  NAND2BXL U203 ( .AN(b[1]), .B(n33), .Y(n127) );
  NAND2XL U204 ( .A(b[2]), .B(n36), .Y(n407) );
  XNOR2X1 U205 ( .A(n141), .B(n174), .Y(n358) );
  XOR2X1 U206 ( .A(n263), .B(n174), .Y(n202) );
  XNOR2X1 U207 ( .A(n67), .B(n4), .Y(n305) );
  XOR2X1 U208 ( .A(n141), .B(n374), .Y(n63) );
  XOR3X2 U209 ( .A(n359), .B(n358), .C(n357), .Y(c[10]) );
  NAND3X1 U210 ( .A(n326), .B(n325), .C(n324), .Y(n381) );
  NAND3X1 U211 ( .A(n52), .B(n319), .C(n321), .Y(n325) );
  XOR2X1 U212 ( .A(n435), .B(n436), .Y(n173) );
  XNOR3X2 U213 ( .A(n63), .B(n175), .C(n196), .Y(n221) );
  NOR2X1 U214 ( .A(n52), .B(n320), .Y(n322) );
  XOR3X2 U215 ( .A(n202), .B(n262), .C(n196), .Y(n203) );
  XNOR3X2 U216 ( .A(n372), .B(n371), .C(n370), .Y(c[11]) );
  XNOR3X2 U217 ( .A(n362), .B(n361), .C(n360), .Y(n372) );
  XOR2X1 U218 ( .A(n367), .B(n366), .Y(n371) );
  XNOR3X2 U219 ( .A(n305), .B(n77), .C(n247), .Y(c[5]) );
  XNOR3X2 U220 ( .A(n456), .B(n246), .C(n240), .Y(n247) );
  XOR2X1 U221 ( .A(n239), .B(n457), .Y(n240) );
  XNOR2X1 U222 ( .A(n459), .B(n458), .Y(n246) );
  XNOR3X2 U223 ( .A(n332), .B(n331), .C(n330), .Y(c[8]) );
  XOR2X1 U224 ( .A(n304), .B(n303), .Y(n332) );
  XNOR2X1 U225 ( .A(n328), .B(n327), .Y(n330) );
  XNOR3X2 U226 ( .A(n314), .B(n306), .C(n305), .Y(n331) );
  INVX1 U227 ( .A(n363), .Y(n374) );
  NOR2X1 U228 ( .A(n382), .B(n384), .Y(n404) );
  XOR3X2 U229 ( .A(n64), .B(n65), .C(n66), .Y(n357) );
  XNOR3X2 U230 ( .A(n395), .B(n394), .C(n393), .Y(n64) );
  XOR2X1 U231 ( .A(n350), .B(n349), .Y(n65) );
  XNOR2X1 U232 ( .A(n356), .B(n355), .Y(n66) );
  XOR2X1 U233 ( .A(n224), .B(n223), .Y(n238) );
  XOR3X2 U234 ( .A(n235), .B(n234), .C(n233), .Y(n236) );
  INVX1 U235 ( .A(n365), .Y(n174) );
  XOR3X2 U236 ( .A(n68), .B(n74), .C(n220), .Y(n67) );
  XNOR2X1 U237 ( .A(n213), .B(n212), .Y(n68) );
  XOR2X1 U238 ( .A(n452), .B(n453), .Y(n74) );
  XOR2X1 U239 ( .A(n381), .B(n5), .Y(n368) );
  XNOR3X2 U240 ( .A(n78), .B(n265), .C(n264), .Y(c[6]) );
  XNOR3X2 U241 ( .A(n374), .B(n263), .C(n262), .Y(n264) );
  XOR2X1 U242 ( .A(n423), .B(n422), .Y(c[12]) );
  XOR2X1 U243 ( .A(n421), .B(n420), .Y(n422) );
  INVX1 U244 ( .A(n323), .Y(n319) );
  INVX1 U245 ( .A(n85), .Y(n180) );
  XNOR2X1 U246 ( .A(n289), .B(n4), .Y(n78) );
  XOR2X1 U247 ( .A(n302), .B(n301), .Y(c[7]) );
  XOR2X1 U248 ( .A(n204), .B(n203), .Y(c[3]) );
  XNOR3X2 U249 ( .A(n222), .B(n266), .C(n221), .Y(c[4]) );
  XNOR3X2 U250 ( .A(n78), .B(n348), .C(n347), .Y(c[9]) );
  NOR2XL U251 ( .A(n480), .B(n382), .Y(n474) );
  OAI21XL U252 ( .A0(n27), .A1(n486), .B0(n10), .Y(n490) );
  OAI21XL U253 ( .A0(n26), .A1(n488), .B0(n8), .Y(n489) );
  OAI21XL U254 ( .A0(n22), .A1(n486), .B0(n10), .Y(n445) );
  OAI21XL U255 ( .A0(n101), .A1(n488), .B0(n8), .Y(n444) );
  OAI21XL U256 ( .A0(n36), .A1(n375), .B0(n10), .Y(n391) );
  OAI21XL U257 ( .A0(n27), .A1(n488), .B0(n8), .Y(n392) );
  AOI22X1 U258 ( .A0(a[4]), .A1(n455), .B0(a[5]), .B1(n454), .Y(n456) );
  OAI21XL U259 ( .A0(a[5]), .A1(n375), .B0(n10), .Y(n455) );
  OAI21XL U260 ( .A0(n102), .A1(n488), .B0(n8), .Y(n454) );
  OAI21XL U261 ( .A0(n104), .A1(n486), .B0(n9), .Y(n464) );
  XNOR3X2 U262 ( .A(n439), .B(n440), .C(n193), .Y(n194) );
  NAND3X1 U263 ( .A(n192), .B(n191), .C(n190), .Y(n195) );
  NAND2X1 U264 ( .A(n24), .B(n30), .Y(n440) );
  OAI21XL U265 ( .A0(n103), .A1(n488), .B0(n487), .Y(n463) );
  OAI21XL U266 ( .A0(n19), .A1(n11), .B0(n8), .Y(n431) );
  OAI21XL U267 ( .A0(n22), .A1(n488), .B0(n8), .Y(n448) );
  OAI21XL U268 ( .A0(a[6]), .A1(n11), .B0(n8), .Y(n472) );
  XNOR3X2 U269 ( .A(n428), .B(n152), .C(n151), .Y(n153) );
  XNOR3X2 U270 ( .A(n148), .B(n147), .C(n146), .Y(n154) );
  INVX1 U271 ( .A(b[2]), .Y(n480) );
  NAND2X1 U272 ( .A(n30), .B(n318), .Y(n321) );
  XOR3X2 U273 ( .A(n179), .B(n178), .C(n177), .Y(n189) );
  NAND2X1 U274 ( .A(b[8]), .B(a[8]), .Y(n178) );
  NAND2X1 U275 ( .A(n96), .B(n105), .Y(n179) );
  XOR2X1 U276 ( .A(n261), .B(n260), .Y(n289) );
  XOR2X1 U277 ( .A(n259), .B(n254), .Y(n260) );
  XNOR3X2 U278 ( .A(n253), .B(n252), .C(n251), .Y(n261) );
  OAI2BB1X1 U279 ( .A0N(n13), .A1N(n126), .B0(n122), .Y(n365) );
  OAI21XL U280 ( .A0(n119), .A1(n377), .B0(n17), .Y(n122) );
  NOR2BX1 U281 ( .AN(a[11]), .B(n86), .Y(n165) );
  XNOR2X1 U282 ( .A(n316), .B(n315), .Y(n323) );
  NAND2X1 U283 ( .A(n35), .B(n98), .Y(n315) );
  XOR2X1 U284 ( .A(n140), .B(n139), .Y(n196) );
  XNOR3X2 U285 ( .A(n386), .B(n138), .C(n137), .Y(n139) );
  XNOR3X2 U286 ( .A(n133), .B(n132), .C(n131), .Y(n140) );
  XNOR3X2 U287 ( .A(n373), .B(n335), .C(n334), .Y(n348) );
  XOR2X1 U288 ( .A(n333), .B(n493), .Y(n334) );
  XNOR2X1 U289 ( .A(n494), .B(n491), .Y(n335) );
  NAND2X1 U290 ( .A(b[4]), .B(n24), .Y(n402) );
  XOR2X1 U291 ( .A(n288), .B(n286), .Y(n300) );
  NAND2X1 U292 ( .A(n100), .B(n12), .Y(n286) );
  XOR2X1 U293 ( .A(n163), .B(n162), .Y(n169) );
  XOR2X1 U294 ( .A(n150), .B(n149), .Y(n152) );
  XOR2X1 U295 ( .A(n388), .B(n389), .Y(n138) );
  NAND2X1 U296 ( .A(n102), .B(n29), .Y(n388) );
  XOR3X2 U297 ( .A(n414), .B(n415), .C(n381), .Y(n423) );
  XOR2X1 U298 ( .A(n411), .B(n410), .Y(n412) );
  XNOR3X2 U299 ( .A(n475), .B(n278), .C(n266), .Y(n302) );
  XOR3X2 U300 ( .A(n476), .B(n477), .C(n474), .Y(n278) );
  AOI22X1 U301 ( .A0(a[6]), .A1(n473), .B0(n24), .B1(n472), .Y(n475) );
  NAND2X1 U302 ( .A(n102), .B(b[3]), .Y(n477) );
  XNOR3X2 U303 ( .A(n63), .B(n443), .C(n176), .Y(n204) );
  NOR2X1 U304 ( .A(n383), .B(n385), .Y(n443) );
  XNOR2X1 U305 ( .A(n446), .B(n447), .Y(n176) );
  INVX1 U306 ( .A(n86), .Y(n385) );
  XOR2X1 U307 ( .A(n409), .B(n408), .Y(n410) );
  XOR2X1 U308 ( .A(n468), .B(n467), .Y(n469) );
  NAND2X1 U309 ( .A(n102), .B(b[4]), .Y(n483) );
  OAI2BB1X1 U310 ( .A0N(n33), .A1N(n214), .B0(n85), .Y(n217) );
  NAND2X1 U311 ( .A(n104), .B(n29), .Y(n435) );
  OAI2BB1X1 U312 ( .A0N(n30), .A1N(n298), .B0(n297), .Y(n299) );
  OAI21XL U313 ( .A0(n296), .A1(n377), .B0(n16), .Y(n297) );
  OAI2BB1X1 U314 ( .A0N(n86), .A1N(n167), .B0(n166), .Y(n168) );
  OAI21XL U315 ( .A0(n165), .A1(n180), .B0(n87), .Y(n166) );
  INVX1 U316 ( .A(n87), .Y(n164) );
  XNOR3X2 U317 ( .A(n80), .B(n81), .C(n387), .Y(n131) );
  XOR3X2 U318 ( .A(n136), .B(n135), .C(n134), .Y(n137) );
  XOR2X1 U319 ( .A(n434), .B(n433), .Y(n438) );
  NOR2X1 U320 ( .A(n383), .B(n480), .Y(n433) );
  AOI22X1 U321 ( .A0(n19), .A1(n432), .B0(n20), .B1(n431), .Y(n434) );
  OAI21XL U322 ( .A0(n20), .A1(n375), .B0(n10), .Y(n432) );
  XNOR3X2 U323 ( .A(n346), .B(n343), .C(n339), .Y(n347) );
  XOR3X2 U324 ( .A(n338), .B(n337), .C(n336), .Y(n339) );
  XOR2X1 U325 ( .A(n381), .B(n492), .Y(n346) );
  AOI21X1 U326 ( .A0(n95), .A1(n217), .B0(n216), .Y(n219) );
  OAI2BB1X1 U327 ( .A0N(n16), .A1N(n250), .B0(n249), .Y(n251) );
  OAI21XL U328 ( .A0(n248), .A1(n377), .B0(n96), .Y(n249) );
  XNOR3X2 U329 ( .A(n390), .B(n358), .C(n196), .Y(c[0]) );
  XOR2X1 U330 ( .A(n466), .B(n465), .Y(n470) );
  AOI22X1 U331 ( .A0(n103), .A1(n464), .B0(n104), .B1(n463), .Y(n466) );
  NAND2X1 U332 ( .A(n92), .B(n24), .Y(n406) );
  XOR2X1 U333 ( .A(n471), .B(n462), .Y(n265) );
  XOR2X1 U334 ( .A(n461), .B(n460), .Y(n462) );
  XOR2X1 U335 ( .A(n470), .B(n469), .Y(n471) );
  NAND2X1 U336 ( .A(n92), .B(a[1]), .Y(n461) );
  OAI21XL U337 ( .A0(n181), .A1(n180), .B0(n92), .Y(n182) );
  OAI21XL U338 ( .A0(n187), .A1(n377), .B0(n87), .Y(n188) );
  OAI21XL U339 ( .A0(n26), .A1(n375), .B0(n10), .Y(n479) );
  OAI21XL U340 ( .A0(n24), .A1(n488), .B0(n8), .Y(n478) );
  OAI21XL U341 ( .A0(n33), .A1(n375), .B0(n10), .Y(n398) );
  OAI21XL U342 ( .A0(n36), .A1(n488), .B0(n8), .Y(n397) );
  XOR2X1 U343 ( .A(n451), .B(n211), .Y(n222) );
  XOR3X2 U344 ( .A(n210), .B(n205), .C(n450), .Y(n211) );
  NOR2X1 U345 ( .A(n480), .B(n485), .Y(n450) );
  NAND2BXL U346 ( .AN(n96), .B(n38), .Y(n226) );
  OAI2BB1X1 U347 ( .A0N(n86), .A1N(n145), .B0(n144), .Y(n147) );
  OAI21XL U348 ( .A0(n143), .A1(n377), .B0(b[2]), .Y(n144) );
  NOR2BX1 U349 ( .AN(a[12]), .B(n86), .Y(n143) );
  AND2X2 U350 ( .A(n99), .B(a[3]), .Y(n155) );
  XNOR3X2 U351 ( .A(n82), .B(n83), .C(n427), .Y(n146) );
  AND2X2 U352 ( .A(n35), .B(n92), .Y(n170) );
  XNOR2X1 U353 ( .A(n429), .B(n426), .Y(n151) );
  XNOR2X1 U354 ( .A(n441), .B(n442), .Y(n193) );
  INVX1 U355 ( .A(n97), .Y(n320) );
  INVX1 U356 ( .A(n92), .Y(n214) );
  OAI21XL U357 ( .A0(n102), .A1(n375), .B0(n10), .Y(n449) );
  OAI21XL U358 ( .A0(n24), .A1(n375), .B0(n10), .Y(n473) );
  NAND2X1 U359 ( .A(n101), .B(n30), .Y(n396) );
  XOR2X1 U360 ( .A(n364), .B(n363), .Y(n84) );
  NAND2X1 U361 ( .A(n100), .B(n31), .Y(n351) );
  NAND2X1 U362 ( .A(n30), .B(a[1]), .Y(n352) );
  XOR2X1 U363 ( .A(n354), .B(n353), .Y(n355) );
  XOR2X1 U364 ( .A(n419), .B(n418), .Y(n420) );
  XOR2X1 U365 ( .A(n484), .B(n481), .Y(n327) );
  AND2X2 U366 ( .A(n86), .B(a[1]), .Y(n205) );
  NAND2X1 U367 ( .A(b[5]), .B(n101), .Y(n288) );
  AND2X2 U368 ( .A(n24), .B(b[2]), .Y(n491) );
  NAND2X1 U369 ( .A(n86), .B(n24), .Y(n395) );
  NAND2X1 U370 ( .A(n100), .B(n30), .Y(n338) );
  NAND2X1 U371 ( .A(a[6]), .B(n92), .Y(n362) );
  INVX1 U372 ( .A(n100), .Y(n383) );
  XOR2X1 U373 ( .A(n417), .B(n416), .Y(n421) );
  AOI22X1 U374 ( .A0(a[0]), .A1(n425), .B0(n19), .B1(n424), .Y(n430) );
  OAI21XL U375 ( .A0(n19), .A1(n375), .B0(n10), .Y(n425) );
  OAI21XL U376 ( .A0(n100), .A1(n11), .B0(n8), .Y(n424) );
  XOR2X1 U377 ( .A(n403), .B(n400), .Y(n369) );
  NOR2X1 U378 ( .A(n399), .B(n480), .Y(n400) );
  INVX1 U379 ( .A(n101), .Y(n485) );
  BUFX3 U380 ( .A(a[4]), .Y(n102) );
  BUFX3 U381 ( .A(a[6]), .Y(n104) );
  BUFX3 U382 ( .A(a[2]), .Y(n101) );
  BUFX3 U383 ( .A(a[5]), .Y(n103) );
  BUFX3 U384 ( .A(b[11]), .Y(n98) );
  BUFX3 U385 ( .A(a[9]), .Y(n105) );
  BUFX3 U386 ( .A(b[10]), .Y(n97) );
  BUFX3 U387 ( .A(b[4]), .Y(n87) );
  BUFX3 U388 ( .A(b[7]), .Y(n96) );
  BUFX3 U389 ( .A(b[3]), .Y(n86) );
  BUFX3 U390 ( .A(b[5]), .Y(n92) );
  BUFX3 U391 ( .A(b[6]), .Y(n95) );
  BUFX3 U392 ( .A(b[12]), .Y(n99) );
  INVX1 U393 ( .A(b[1]), .Y(n375) );
  XOR2X1 U394 ( .A(n380), .B(n407), .Y(n411) );
  OAI2BB1X1 U395 ( .A0N(b[2]), .A1N(n130), .B0(n129), .Y(n132) );
  OAI21XL U396 ( .A0(n128), .A1(n377), .B0(b[1]), .Y(n129) );
  NOR2BX1 U397 ( .AN(n38), .B(b[2]), .Y(n128) );
  BUFX3 U398 ( .A(a[0]), .Y(n100) );
  AOI21XL U399 ( .A0(n317), .A1(n226), .B0(n225), .Y(n230) );
  AOI21XL U400 ( .A0(n317), .A1(n215), .B0(n214), .Y(n216) );
  OAI2BB1XL U401 ( .A0N(a[12]), .A1N(n164), .B0(n317), .Y(n167) );
  XOR2X4 U402 ( .A(n110), .B(n109), .Y(n373) );
endmodule


module multiplier_4 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n36, n37, n38, n39, n47, n49, n50, n51, n52, n53,
         n54, n55, n57, n58, n59, n61, n63, n64, n74, n77, n81, n83, n84, n85,
         n86, n87, n92, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n122, n127, n128, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n202, n203, n204, n205, n210,
         n211, n212, n213, n214, n215, n216, n217, n219, n220, n221, n239,
         n240, n246, n247, n248, n249, n250, n251, n252, n253, n254, n259,
         n260, n261, n262, n263, n264, n265, n266, n286, n288, n289, n290,
         n291, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n311, n314, n315, n316, n317, n318, n319, n320, n321, n323,
         n324, n325, n326, n327, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542;

  OAI2BB1XL U1 ( .A0N(n15), .A1N(n39), .B0(n370), .Y(n303) );
  CLKINVXL U2 ( .A(n370), .Y(n317) );
  AOI21XL U3 ( .A0(n370), .A1(n260), .B0(n395), .Y(n261) );
  BUFX4 U4 ( .A(a[12]), .Y(n100) );
  OAI21XL U5 ( .A0(n1), .A1(n85), .B0(n370), .Y(n239) );
  INVX1 U6 ( .A(n39), .Y(n1) );
  OAI221XL U7 ( .A0(n106), .A1(n57), .B0(n5), .B1(n375), .C0(n371), .Y(n372)
         );
  AND2X2 U8 ( .A(n74), .B(n99), .Y(n523) );
  NOR2X1 U9 ( .A(n33), .B(n9), .Y(n306) );
  NOR2X1 U10 ( .A(n19), .B(n375), .Y(n301) );
  NAND2BX1 U11 ( .AN(n167), .B(n169), .Y(n170) );
  OAI21XL U12 ( .A0(n2), .A1(n74), .B0(n370), .Y(n142) );
  INVX1 U13 ( .A(n38), .Y(n2) );
  NOR2BX1 U14 ( .AN(n39), .B(n100), .Y(n373) );
  OR2X2 U15 ( .A(n168), .B(n165), .Y(n174) );
  AOI22XL U16 ( .A0(a[10]), .A1(n405), .B0(n32), .B1(n404), .Y(n407) );
  NOR2X1 U17 ( .A(n375), .B(n77), .Y(n140) );
  XOR2X1 U18 ( .A(n298), .B(n3), .Y(n337) );
  OAI21XL U19 ( .A0(n375), .A1(b[10]), .B0(n316), .Y(n320) );
  NAND3X1 U20 ( .A(n168), .B(n165), .C(n167), .Y(n173) );
  NOR2X1 U21 ( .A(n522), .B(n30), .Y(n415) );
  XOR3X2 U22 ( .A(n353), .B(n337), .C(n352), .Y(c[10]) );
  XNOR3X2 U23 ( .A(n381), .B(n469), .C(n180), .Y(c[2]) );
  OAI2BB1X2 U24 ( .A0N(n39), .A1N(n9), .B0(n370), .Y(n103) );
  AOI21X1 U25 ( .A0(n316), .A1(n101), .B0(n9), .Y(n102) );
  INVX1 U26 ( .A(n213), .Y(n219) );
  XNOR2X2 U27 ( .A(n105), .B(n104), .Y(n139) );
  NAND2BX2 U28 ( .AN(n100), .B(n38), .Y(n370) );
  INVX1 U29 ( .A(n21), .Y(n22) );
  NAND2BX1 U30 ( .AN(a[11]), .B(n100), .Y(n316) );
  INVX2 U31 ( .A(n139), .Y(n333) );
  BUFX3 U32 ( .A(a[11]), .Y(n39) );
  XNOR3X2 U33 ( .A(n306), .B(n305), .C(n304), .Y(n3) );
  INVX1 U34 ( .A(b[0]), .Y(n4) );
  NAND2X1 U35 ( .A(b[0]), .B(n534), .Y(n5) );
  NAND2X1 U36 ( .A(b[0]), .B(n534), .Y(n55) );
  BUFX3 U37 ( .A(n57), .Y(n6) );
  NAND2X1 U38 ( .A(b[1]), .B(n535), .Y(n57) );
  INVX1 U39 ( .A(n395), .Y(n7) );
  INVX1 U40 ( .A(n396), .Y(n8) );
  BUFX3 U41 ( .A(b[3]), .Y(n77) );
  INVX1 U42 ( .A(b[10]), .Y(n9) );
  INVXL U43 ( .A(n9), .Y(n10) );
  INVX1 U44 ( .A(n190), .Y(n11) );
  INVX1 U45 ( .A(n394), .Y(n12) );
  INVX1 U46 ( .A(n387), .Y(n13) );
  INVX1 U47 ( .A(n254), .Y(n14) );
  INVX1 U48 ( .A(b[8]), .Y(n15) );
  INVX1 U49 ( .A(n15), .Y(n16) );
  INVX1 U50 ( .A(n15), .Y(n17) );
  INVX1 U51 ( .A(b[9]), .Y(n18) );
  INVX1 U52 ( .A(n18), .Y(n19) );
  INVX1 U53 ( .A(n18), .Y(n20) );
  INVX1 U54 ( .A(b[11]), .Y(n21) );
  INVX1 U55 ( .A(n533), .Y(n23) );
  INVX1 U56 ( .A(n466), .Y(n24) );
  INVX1 U57 ( .A(n502), .Y(n25) );
  INVX1 U58 ( .A(a[7]), .Y(n26) );
  INVXL U59 ( .A(n26), .Y(n27) );
  INVX1 U60 ( .A(a[8]), .Y(n28) );
  INVX1 U61 ( .A(n28), .Y(n29) );
  INVX1 U62 ( .A(a[9]), .Y(n30) );
  INVX1 U63 ( .A(n30), .Y(n31) );
  INVX1 U64 ( .A(n30), .Y(n32) );
  INVX1 U65 ( .A(a[10]), .Y(n33) );
  INVX1 U66 ( .A(n33), .Y(n34) );
  INVXL U67 ( .A(n33), .Y(n36) );
  AND2X2 U68 ( .A(n34), .B(n86), .Y(n104) );
  INVX1 U69 ( .A(n375), .Y(n37) );
  OAI21X1 U70 ( .A0(n378), .A1(n377), .B0(n376), .Y(n452) );
  INVX2 U71 ( .A(n496), .Y(n385) );
  XOR2X2 U72 ( .A(n468), .B(n467), .Y(n496) );
  XOR3X4 U73 ( .A(n385), .B(n384), .C(n383), .Y(n494) );
  AOI21X2 U74 ( .A0(b[11]), .A1(n103), .B0(n102), .Y(n105) );
  BUFX3 U75 ( .A(b[4]), .Y(n81) );
  BUFX2 U76 ( .A(a[11]), .Y(n38) );
  OAI2BB1XL U77 ( .A0N(n39), .A1N(n81), .B0(n396), .Y(n376) );
  NOR2BX1 U78 ( .AN(n38), .B(n81), .Y(n166) );
  XOR2X1 U79 ( .A(n495), .B(n494), .Y(c[5]) );
  XNOR3X2 U80 ( .A(n367), .B(n366), .C(n365), .Y(c[11]) );
  NOR2BX1 U81 ( .AN(n38), .B(n20), .Y(n318) );
  NAND2XL U82 ( .A(n96), .B(n22), .Y(n146) );
  INVX1 U83 ( .A(n83), .Y(n190) );
  AOI21X1 U84 ( .A0(n84), .A1(n193), .B0(n192), .Y(n212) );
  NAND2X1 U85 ( .A(n85), .B(n31), .Y(n163) );
  NAND2X1 U86 ( .A(n16), .B(a[8]), .Y(n162) );
  NAND2XL U87 ( .A(n96), .B(n77), .Y(n506) );
  NAND2XL U88 ( .A(n8), .B(n29), .Y(n418) );
  NAND2XL U89 ( .A(n97), .B(n77), .Y(n515) );
  NAND2XL U90 ( .A(a[8]), .B(n83), .Y(n63) );
  NAND2XL U91 ( .A(n77), .B(a[6]), .Y(n541) );
  AND2X1 U92 ( .A(n29), .B(n74), .Y(n406) );
  INVXL U93 ( .A(n368), .Y(n179) );
  XOR3X2 U94 ( .A(n49), .B(n286), .C(n266), .Y(n47) );
  XNOR2X1 U95 ( .A(n253), .B(n252), .Y(n49) );
  NOR2XL U96 ( .A(n387), .B(n395), .Y(n419) );
  NOR2XL U97 ( .A(n389), .B(n396), .Y(n474) );
  NOR2XL U98 ( .A(n388), .B(n395), .Y(n516) );
  XOR3X2 U99 ( .A(n50), .B(n406), .C(n51), .Y(n352) );
  XOR3X2 U100 ( .A(n407), .B(n339), .C(n338), .Y(n50) );
  XNOR3X2 U101 ( .A(n351), .B(n350), .C(n349), .Y(n51) );
  XOR2X1 U102 ( .A(n152), .B(n447), .Y(c[1]) );
  INVXL U103 ( .A(n100), .Y(n375) );
  NAND2XL U104 ( .A(n97), .B(n10), .Y(n445) );
  INVXL U105 ( .A(n38), .Y(n106) );
  AOI22XL U106 ( .A0(n12), .A1(n108), .B0(n22), .B1(n107), .Y(n382) );
  NAND2XL U107 ( .A(n7), .B(n96), .Y(n339) );
  NAND2XL U108 ( .A(n20), .B(n36), .Y(n246) );
  NAND2XL U109 ( .A(n99), .B(n86), .Y(n264) );
  NAND2XL U110 ( .A(n85), .B(n29), .Y(n454) );
  AOI22XL U111 ( .A0(n29), .A1(n537), .B0(n32), .B1(n536), .Y(n539) );
  NAND2XL U112 ( .A(n97), .B(n19), .Y(n401) );
  NAND2XL U113 ( .A(n98), .B(n16), .Y(n402) );
  NAND2XL U114 ( .A(n86), .B(n95), .Y(n147) );
  NAND2BXL U115 ( .AN(n84), .B(n100), .Y(n191) );
  INVXL U116 ( .A(n85), .Y(n395) );
  NAND2XL U117 ( .A(n27), .B(n12), .Y(n249) );
  NAND2XL U118 ( .A(n37), .B(n86), .Y(n216) );
  NAND2XL U119 ( .A(n29), .B(n10), .Y(n263) );
  OAI21XL U120 ( .A0(n318), .A1(n317), .B0(n10), .Y(n319) );
  XNOR3X2 U121 ( .A(n52), .B(n412), .C(n321), .Y(n542) );
  NAND2XL U122 ( .A(n32), .B(n86), .Y(n52) );
  NAND2XL U123 ( .A(a[7]), .B(n20), .Y(n471) );
  OAI2BB1X1 U124 ( .A0N(n77), .A1N(n142), .B0(n141), .Y(n144) );
  NAND2XL U125 ( .A(b[4]), .B(n98), .Y(n540) );
  XNOR3X2 U126 ( .A(n334), .B(n333), .C(n539), .Y(n335) );
  NAND2XL U127 ( .A(n87), .B(n20), .Y(n331) );
  NAND2XL U128 ( .A(n85), .B(n95), .Y(n330) );
  NAND2XL U129 ( .A(n96), .B(b[4]), .Y(n514) );
  NAND2XL U130 ( .A(n36), .B(n77), .Y(n136) );
  NAND2XL U131 ( .A(n99), .B(n10), .Y(n470) );
  NAND2XL U132 ( .A(n74), .B(n36), .Y(n423) );
  NAND2XL U133 ( .A(n84), .B(a[6]), .Y(n420) );
  NAND2XL U134 ( .A(n77), .B(n27), .Y(n409) );
  NAND2XL U135 ( .A(b[4]), .B(n99), .Y(n408) );
  NAND2XL U136 ( .A(b[4]), .B(n29), .Y(n424) );
  NAND2XL U137 ( .A(n99), .B(n19), .Y(n458) );
  NAND2XL U138 ( .A(n17), .B(n92), .Y(n323) );
  NAND2XL U139 ( .A(n87), .B(n7), .Y(n296) );
  NAND2XL U140 ( .A(n14), .B(n87), .Y(n497) );
  NAND2XL U141 ( .A(n97), .B(n81), .Y(n525) );
  NAND2XL U142 ( .A(n31), .B(b[11]), .Y(n299) );
  XOR2X1 U143 ( .A(n205), .B(n204), .Y(n210) );
  NAND2XL U144 ( .A(n83), .B(n36), .Y(n453) );
  NAND2XL U145 ( .A(a[8]), .B(n86), .Y(n300) );
  NAND2XL U146 ( .A(n83), .B(n92), .Y(n498) );
  NAND2XL U147 ( .A(a[7]), .B(n10), .Y(n485) );
  NAND2XL U148 ( .A(n98), .B(n10), .Y(n461) );
  NAND2XL U149 ( .A(n97), .B(n14), .Y(n346) );
  NAND2XL U150 ( .A(n87), .B(n10), .Y(n347) );
  NAND2XL U151 ( .A(n20), .B(n92), .Y(n348) );
  NAND2XL U152 ( .A(n85), .B(n27), .Y(n444) );
  NAND2XL U153 ( .A(n84), .B(a[7]), .Y(n400) );
  NAND2XL U154 ( .A(n13), .B(n11), .Y(n338) );
  NAND2XL U155 ( .A(n84), .B(n34), .Y(n153) );
  NAND2BXL U156 ( .AN(b[11]), .B(n100), .Y(n101) );
  NAND2XL U157 ( .A(a[7]), .B(n17), .Y(n459) );
  NAND2XL U158 ( .A(n95), .B(b[4]), .Y(n505) );
  NAND2XL U159 ( .A(n24), .B(n83), .Y(n518) );
  NAND2XL U160 ( .A(n14), .B(n95), .Y(n517) );
  NAND2XL U161 ( .A(n85), .B(n34), .Y(n195) );
  NAND2XL U162 ( .A(n16), .B(n31), .Y(n194) );
  AOI22XL U163 ( .A0(n36), .A1(n414), .B0(n39), .B1(n413), .Y(n416) );
  NAND2XL U164 ( .A(n84), .B(n96), .Y(n324) );
  XNOR3X2 U165 ( .A(n382), .B(n53), .C(n381), .Y(n383) );
  NAND2XL U166 ( .A(n11), .B(n87), .Y(n53) );
  NAND2XL U167 ( .A(n85), .B(n99), .Y(n399) );
  XOR3X2 U168 ( .A(n54), .B(n311), .C(n337), .Y(n314) );
  NAND2XL U169 ( .A(n14), .B(n92), .Y(n54) );
  OAI2BB1XL U170 ( .A0N(n38), .A1N(n190), .B0(n370), .Y(n193) );
  AOI22XL U171 ( .A0(a[6]), .A1(n511), .B0(n27), .B1(n510), .Y(n513) );
  NAND2XL U172 ( .A(n84), .B(a[8]), .Y(n59) );
  NAND2XL U173 ( .A(n32), .B(n83), .Y(n61) );
  NAND2XL U174 ( .A(n86), .B(n92), .Y(n109) );
  NAND2XL U175 ( .A(b[11]), .B(n95), .Y(n110) );
  NAND2XL U176 ( .A(b[10]), .B(n96), .Y(n111) );
  NAND2XL U177 ( .A(n31), .B(n81), .Y(n64) );
  AOI22XL U178 ( .A0(n27), .A1(n521), .B0(n29), .B1(n520), .Y(n524) );
  NAND2XL U179 ( .A(n83), .B(n27), .Y(n421) );
  NAND2XL U180 ( .A(n87), .B(n12), .Y(n430) );
  NAND2XL U181 ( .A(n77), .B(n32), .Y(n425) );
  NAND2XL U182 ( .A(n22), .B(n36), .Y(n412) );
  NAND2XL U183 ( .A(n97), .B(n86), .Y(n472) );
  NAND2XL U184 ( .A(n98), .B(n22), .Y(n473) );
  NAND2XL U185 ( .A(n98), .B(n20), .Y(n446) );
  NAND2XL U186 ( .A(n99), .B(n17), .Y(n443) );
  INVXL U187 ( .A(n84), .Y(n254) );
  INVXL U188 ( .A(n86), .Y(n394) );
  AND2X1 U189 ( .A(n32), .B(b[10]), .Y(n247) );
  AND2X1 U190 ( .A(n36), .B(n81), .Y(n145) );
  AND2X1 U191 ( .A(n87), .B(b[4]), .Y(n188) );
  AND2X1 U192 ( .A(n97), .B(n83), .Y(n325) );
  OAI21XL U193 ( .A0(n164), .A1(n377), .B0(n81), .Y(n165) );
  AND2X1 U194 ( .A(n27), .B(n74), .Y(n538) );
  XOR2X1 U195 ( .A(n457), .B(n456), .Y(n465) );
  XOR2X1 U196 ( .A(n455), .B(n454), .Y(n456) );
  NAND2XL U197 ( .A(n84), .B(n32), .Y(n455) );
  NAND2XL U198 ( .A(n98), .B(n86), .Y(n203) );
  NAND2XL U199 ( .A(n19), .B(a[8]), .Y(n202) );
  OAI21XL U200 ( .A0(n166), .A1(n373), .B0(n83), .Y(n167) );
  INVX2 U201 ( .A(n77), .Y(n396) );
  NAND2XL U202 ( .A(n17), .B(n95), .Y(n350) );
  NAND2XL U203 ( .A(n87), .B(n22), .Y(n361) );
  NAND2XL U204 ( .A(a[6]), .B(n11), .Y(n356) );
  NAND2XL U205 ( .A(n13), .B(n14), .Y(n357) );
  NAND2XL U206 ( .A(n25), .B(n7), .Y(n358) );
  NAND2XL U207 ( .A(n81), .B(n27), .Y(n417) );
  NAND2XL U208 ( .A(n24), .B(n20), .Y(n433) );
  NAND2XL U209 ( .A(n24), .B(n17), .Y(n411) );
  NAND2XL U210 ( .A(n81), .B(a[1]), .Y(n490) );
  NAND2XL U211 ( .A(n92), .B(n22), .Y(n435) );
  NAND2XL U212 ( .A(n23), .B(n20), .Y(n410) );
  AND2X1 U213 ( .A(n17), .B(a[0]), .Y(n531) );
  NAND2XL U214 ( .A(n98), .B(n8), .Y(n526) );
  NAND2XL U215 ( .A(n23), .B(n10), .Y(n436) );
  NAND2XL U216 ( .A(a[1]), .B(n10), .Y(n360) );
  NAND2XL U217 ( .A(n25), .B(n17), .Y(n434) );
  NAND2XL U218 ( .A(n370), .B(n128), .Y(n133) );
  NAND2BXL U219 ( .AN(b[1]), .B(n39), .Y(n128) );
  AOI2BB2XL U220 ( .B0(b[0]), .B1(n377), .A0N(n370), .A1N(n369), .Y(n371) );
  INVXL U221 ( .A(b[1]), .Y(n369) );
  XNOR2X1 U222 ( .A(n333), .B(n359), .Y(n368) );
  XOR2X1 U223 ( .A(n58), .B(n385), .Y(n288) );
  INVX1 U224 ( .A(n214), .Y(n152) );
  INVX1 U225 ( .A(n316), .Y(n377) );
  XOR2X1 U226 ( .A(n542), .B(n3), .Y(n355) );
  XOR2X1 U227 ( .A(n213), .B(n380), .Y(n290) );
  XNOR3X2 U228 ( .A(n179), .B(n178), .C(n381), .Y(n214) );
  XOR3X2 U229 ( .A(n265), .B(n264), .C(n263), .Y(n266) );
  XNOR3X2 U230 ( .A(n179), .B(n219), .C(n178), .Y(n181) );
  XNOR2X1 U231 ( .A(n496), .B(n382), .Y(n180) );
  NOR2X1 U232 ( .A(n373), .B(n396), .Y(n374) );
  XOR3X2 U233 ( .A(n516), .B(n47), .C(n386), .Y(n397) );
  XNOR3X2 U234 ( .A(n219), .B(n509), .C(n217), .Y(n289) );
  XOR2X1 U235 ( .A(n216), .B(n499), .Y(n217) );
  XOR2X1 U236 ( .A(n508), .B(n507), .Y(n509) );
  XOR2X1 U237 ( .A(n498), .B(n497), .Y(n499) );
  XOR3X2 U238 ( .A(n364), .B(n363), .C(n362), .Y(n365) );
  XOR2X1 U239 ( .A(n410), .B(n411), .Y(n363) );
  XNOR3X2 U240 ( .A(n417), .B(n361), .C(n360), .Y(n362) );
  XOR2X1 U241 ( .A(n382), .B(n359), .Y(n364) );
  INVX1 U242 ( .A(n216), .Y(n359) );
  INVX1 U243 ( .A(n386), .Y(n380) );
  XOR2X1 U244 ( .A(n289), .B(n288), .Y(c[6]) );
  XOR2X1 U245 ( .A(n440), .B(n439), .Y(c[12]) );
  XNOR2X1 U246 ( .A(n298), .B(n47), .Y(n58) );
  XOR2X1 U247 ( .A(n530), .B(n529), .Y(n532) );
  XOR2X1 U248 ( .A(n528), .B(n527), .Y(n529) );
  XOR2X1 U249 ( .A(n397), .B(n519), .Y(n530) );
  XOR2X1 U250 ( .A(n526), .B(n525), .Y(n527) );
  INVX1 U251 ( .A(n168), .Y(n169) );
  XOR2X1 U252 ( .A(n479), .B(n474), .Y(n182) );
  XOR2X1 U253 ( .A(n478), .B(n477), .Y(n479) );
  NOR2X1 U254 ( .A(n388), .B(n522), .Y(n477) );
  XOR3X2 U255 ( .A(n355), .B(n531), .C(n532), .Y(c[8]) );
  XOR2X1 U256 ( .A(n315), .B(n314), .Y(c[7]) );
  XNOR3X2 U257 ( .A(n182), .B(n181), .C(n180), .Y(c[3]) );
  XNOR3X2 U258 ( .A(n215), .B(n290), .C(n214), .Y(c[4]) );
  XNOR3X2 U259 ( .A(n336), .B(n58), .C(n335), .Y(c[9]) );
  NOR2X1 U260 ( .A(n522), .B(n387), .Y(n512) );
  OAI21XL U261 ( .A0(n22), .A1(n106), .B0(n370), .Y(n108) );
  OAI21XL U262 ( .A0(n32), .A1(n369), .B0(n6), .Y(n537) );
  OAI21XL U263 ( .A0(n29), .A1(n4), .B0(n55), .Y(n536) );
  AOI22X1 U264 ( .A0(n95), .A1(n476), .B0(n96), .B1(n475), .Y(n478) );
  OAI21XL U265 ( .A0(n96), .A1(n369), .B0(n57), .Y(n476) );
  OAI21XL U266 ( .A0(n95), .A1(n4), .B0(n55), .Y(n475) );
  OAI21XL U267 ( .A0(n36), .A1(n369), .B0(n57), .Y(n404) );
  OAI21XL U268 ( .A0(n32), .A1(n4), .B0(n55), .Y(n405) );
  NOR2X1 U269 ( .A(n262), .B(n261), .Y(n286) );
  NAND2BX1 U270 ( .AN(n84), .B(n38), .Y(n260) );
  OAI2BB1X1 U271 ( .A0N(n20), .A1N(n320), .B0(n319), .Y(n321) );
  OAI21XL U272 ( .A0(n99), .A1(n369), .B0(n57), .Y(n501) );
  OAI21XL U273 ( .A0(n29), .A1(n369), .B0(n57), .Y(n521) );
  OAI21XL U274 ( .A0(n97), .A1(n369), .B0(n57), .Y(n481) );
  OAI21XL U275 ( .A0(n27), .A1(n534), .B0(n57), .Y(n511) );
  OAI21XL U276 ( .A0(n38), .A1(n369), .B0(n57), .Y(n414) );
  OAI21XL U277 ( .A0(n98), .A1(n4), .B0(n55), .Y(n500) );
  OAI21XL U278 ( .A0(n27), .A1(n4), .B0(n5), .Y(n520) );
  OAI21XL U279 ( .A0(n92), .A1(n535), .B0(n55), .Y(n448) );
  OAI21XL U280 ( .A0(n96), .A1(n4), .B0(n55), .Y(n480) );
  AOI22X1 U281 ( .A0(n25), .A1(n487), .B0(n13), .B1(n486), .Y(n488) );
  OAI21XL U282 ( .A0(n13), .A1(n369), .B0(n6), .Y(n487) );
  OAI21XL U283 ( .A0(n25), .A1(n535), .B0(n5), .Y(n486) );
  OAI21XL U284 ( .A0(a[6]), .A1(n4), .B0(n5), .Y(n510) );
  OAI21XL U285 ( .A0(n36), .A1(n4), .B0(n5), .Y(n413) );
  INVX1 U286 ( .A(n74), .Y(n522) );
  MXI2X1 U287 ( .A(n375), .B(n374), .S0(n81), .Y(n378) );
  XOR2X1 U288 ( .A(n151), .B(n150), .Y(n381) );
  XNOR3X2 U289 ( .A(n445), .B(n149), .C(n148), .Y(n150) );
  XNOR3X2 U290 ( .A(n145), .B(n144), .C(n143), .Y(n151) );
  XOR2X1 U291 ( .A(n138), .B(n137), .Y(n178) );
  XNOR3X2 U292 ( .A(n399), .B(n127), .C(n122), .Y(n138) );
  XNOR3X2 U293 ( .A(n136), .B(n135), .C(n134), .Y(n137) );
  XOR3X2 U294 ( .A(n163), .B(n162), .C(n153), .Y(n168) );
  XNOR3X2 U295 ( .A(n212), .B(n211), .C(n210), .Y(n386) );
  XNOR2X1 U296 ( .A(n485), .B(n484), .Y(n211) );
  XOR2X1 U297 ( .A(n177), .B(n176), .Y(n213) );
  XNOR3X2 U298 ( .A(n470), .B(n471), .C(n175), .Y(n176) );
  NAND3X1 U299 ( .A(n174), .B(n173), .C(n170), .Y(n177) );
  XOR2X1 U300 ( .A(n251), .B(n250), .Y(n298) );
  XOR2X1 U301 ( .A(n249), .B(n248), .Y(n250) );
  XNOR3X2 U302 ( .A(n247), .B(n246), .C(n240), .Y(n251) );
  NOR2X1 U303 ( .A(n394), .B(n466), .Y(n467) );
  XOR2X1 U304 ( .A(n465), .B(n464), .Y(n468) );
  INVX1 U305 ( .A(n96), .Y(n466) );
  NOR2BX1 U306 ( .AN(n100), .B(n17), .Y(n220) );
  NOR2BX1 U307 ( .AN(n100), .B(n74), .Y(n131) );
  OAI21XL U308 ( .A0(n140), .A1(n377), .B0(n74), .Y(n141) );
  NAND2X1 U309 ( .A(n97), .B(n22), .Y(n460) );
  NAND2X1 U310 ( .A(a[7]), .B(b[11]), .Y(n252) );
  NAND2X1 U311 ( .A(n29), .B(n22), .Y(n248) );
  NAND2X1 U312 ( .A(n99), .B(n22), .Y(n484) );
  XNOR2X1 U313 ( .A(n195), .B(n194), .Y(n205) );
  XOR2X1 U314 ( .A(n506), .B(n505), .Y(n507) );
  XOR2X1 U315 ( .A(n380), .B(n47), .Y(n384) );
  XOR2X1 U316 ( .A(n297), .B(n296), .Y(n311) );
  NAND2X1 U317 ( .A(n11), .B(n95), .Y(n297) );
  XOR2X1 U318 ( .A(n451), .B(n450), .Y(n469) );
  NOR2X1 U319 ( .A(n389), .B(n522), .Y(n450) );
  AOI22X1 U320 ( .A0(n92), .A1(n449), .B0(n23), .B1(n448), .Y(n451) );
  OAI21XL U321 ( .A0(n23), .A1(n369), .B0(n57), .Y(n449) );
  XOR2X1 U322 ( .A(n147), .B(n146), .Y(n149) );
  XOR2X1 U323 ( .A(n401), .B(n402), .Y(n127) );
  XNOR3X2 U324 ( .A(n513), .B(n291), .C(n290), .Y(n315) );
  XOR3X2 U325 ( .A(n514), .B(n515), .C(n512), .Y(n291) );
  XOR2X1 U326 ( .A(n203), .B(n202), .Y(n204) );
  XOR2X1 U327 ( .A(n463), .B(n462), .Y(n464) );
  XOR2X1 U328 ( .A(n459), .B(n458), .Y(n463) );
  XOR2X1 U329 ( .A(n461), .B(n460), .Y(n462) );
  XOR2X1 U330 ( .A(n427), .B(n426), .Y(n428) );
  XOR2X1 U331 ( .A(n425), .B(n424), .Y(n426) );
  XOR2X1 U332 ( .A(n372), .B(n423), .Y(n427) );
  NAND2X1 U333 ( .A(n16), .B(n34), .Y(n253) );
  XNOR3X2 U334 ( .A(n416), .B(n355), .C(n354), .Y(n367) );
  XNOR2X1 U335 ( .A(n415), .B(n418), .Y(n354) );
  XNOR3X2 U336 ( .A(n327), .B(n326), .C(n542), .Y(n336) );
  XOR2X1 U337 ( .A(n324), .B(n323), .Y(n327) );
  XOR2X1 U338 ( .A(n538), .B(n325), .Y(n326) );
  OAI2BB1X1 U339 ( .A0N(n20), .A1N(n303), .B0(n302), .Y(n304) );
  OAI21XL U340 ( .A0(n301), .A1(n377), .B0(n17), .Y(n302) );
  XNOR3X2 U341 ( .A(n59), .B(n61), .C(n444), .Y(n143) );
  XNOR3X2 U342 ( .A(n63), .B(n64), .C(n400), .Y(n134) );
  XOR3X2 U343 ( .A(n540), .B(n541), .C(n332), .Y(n334) );
  XOR2X1 U344 ( .A(n300), .B(n299), .Y(n305) );
  XNOR3X2 U345 ( .A(n111), .B(n110), .C(n109), .Y(n122) );
  NAND2X1 U346 ( .A(n19), .B(n31), .Y(n265) );
  OAI2BB1X1 U347 ( .A0N(n17), .A1N(n239), .B0(n221), .Y(n240) );
  OAI21XL U348 ( .A0(n220), .A1(n377), .B0(n85), .Y(n221) );
  XNOR3X2 U349 ( .A(n403), .B(n353), .C(n178), .Y(c[0]) );
  XOR2X1 U350 ( .A(n504), .B(n503), .Y(n508) );
  NOR2X1 U351 ( .A(n522), .B(n502), .Y(n503) );
  AOI22X1 U352 ( .A0(n98), .A1(n501), .B0(n99), .B1(n500), .Y(n504) );
  INVX1 U353 ( .A(n97), .Y(n502) );
  XOR2X1 U354 ( .A(n524), .B(n523), .Y(n528) );
  XOR2X1 U355 ( .A(n432), .B(n431), .Y(n440) );
  XNOR2X1 U356 ( .A(n430), .B(n542), .Y(n431) );
  XOR2X1 U357 ( .A(n429), .B(n428), .Y(n432) );
  XOR2X1 U358 ( .A(n453), .B(n452), .Y(n457) );
  XOR2X1 U359 ( .A(n398), .B(n422), .Y(n429) );
  XOR2X1 U360 ( .A(n421), .B(n420), .Y(n422) );
  XOR2X1 U361 ( .A(n368), .B(n419), .Y(n398) );
  XOR2X1 U362 ( .A(n493), .B(n492), .Y(n495) );
  XOR2X1 U363 ( .A(n491), .B(n490), .Y(n492) );
  XOR2X1 U364 ( .A(n489), .B(n488), .Y(n493) );
  NAND2X1 U365 ( .A(n23), .B(n8), .Y(n491) );
  NOR2BX1 U366 ( .AN(n100), .B(n83), .Y(n164) );
  NAND2BX1 U367 ( .AN(n85), .B(n100), .Y(n259) );
  XOR2X1 U368 ( .A(n483), .B(n189), .Y(n215) );
  XOR3X2 U369 ( .A(n188), .B(n187), .C(n482), .Y(n189) );
  AOI22X1 U370 ( .A0(n24), .A1(n481), .B0(n25), .B1(n480), .Y(n483) );
  NOR2X1 U371 ( .A(n522), .B(n533), .Y(n482) );
  INVX1 U372 ( .A(n98), .Y(n387) );
  XNOR2X1 U373 ( .A(n472), .B(n473), .Y(n175) );
  XNOR2X1 U374 ( .A(n446), .B(n443), .Y(n148) );
  AOI22X1 U375 ( .A0(a[0]), .A1(n442), .B0(a[1]), .B1(n441), .Y(n447) );
  OAI21XL U376 ( .A0(a[1]), .A1(n534), .B0(n6), .Y(n442) );
  OAI21XL U377 ( .A0(n87), .A1(n4), .B0(n5), .Y(n441) );
  NOR2X1 U378 ( .A(n389), .B(n4), .Y(n403) );
  XOR2X1 U379 ( .A(n518), .B(n517), .Y(n519) );
  XOR2X1 U380 ( .A(n438), .B(n437), .Y(n439) );
  XOR2X1 U381 ( .A(n434), .B(n433), .Y(n438) );
  XOR2X1 U382 ( .A(n436), .B(n435), .Y(n437) );
  AND2X2 U383 ( .A(n77), .B(n92), .Y(n187) );
  NAND2X1 U384 ( .A(n24), .B(n74), .Y(n489) );
  XOR3X2 U385 ( .A(n348), .B(n347), .C(n346), .Y(n349) );
  XNOR3X2 U386 ( .A(n358), .B(n357), .C(n356), .Y(n366) );
  INVX1 U387 ( .A(n87), .Y(n389) );
  XOR2X1 U388 ( .A(n331), .B(n330), .Y(n332) );
  XOR2X1 U389 ( .A(n409), .B(n408), .Y(n351) );
  INVX1 U390 ( .A(n92), .Y(n388) );
  INVX1 U391 ( .A(n95), .Y(n533) );
  OAI2BB1X1 U392 ( .A0N(n74), .A1N(n133), .B0(n132), .Y(n135) );
  OAI21XL U393 ( .A0(n131), .A1(n377), .B0(b[1]), .Y(n132) );
  BUFX3 U394 ( .A(a[3]), .Y(n96) );
  BUFX3 U395 ( .A(a[6]), .Y(n99) );
  BUFX3 U396 ( .A(a[2]), .Y(n95) );
  BUFX3 U397 ( .A(a[4]), .Y(n97) );
  BUFX3 U398 ( .A(a[5]), .Y(n98) );
  BUFX3 U399 ( .A(b[6]), .Y(n84) );
  BUFX3 U400 ( .A(a[1]), .Y(n92) );
  BUFX3 U401 ( .A(b[12]), .Y(n86) );
  BUFX3 U402 ( .A(b[7]), .Y(n85) );
  BUFX3 U403 ( .A(b[5]), .Y(n83) );
  INVX1 U404 ( .A(b[0]), .Y(n535) );
  INVX1 U405 ( .A(b[1]), .Y(n534) );
  BUFX3 U406 ( .A(b[2]), .Y(n74) );
  BUFX3 U407 ( .A(a[0]), .Y(n87) );
  OAI21XL U408 ( .A0(n12), .A1(n375), .B0(n316), .Y(n107) );
  AOI21X1 U409 ( .A0(n316), .A1(n191), .B0(n190), .Y(n192) );
  AOI21X1 U410 ( .A0(n316), .A1(n259), .B0(n254), .Y(n262) );
  XOR2X1 U411 ( .A(n139), .B(n382), .Y(n353) );
endmodule


module multiplier_3 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n47, n49, n50, n51, n52,
         n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n74, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n92,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n122, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n202,
         n203, n204, n205, n210, n211, n212, n213, n214, n215, n216, n217,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n230,
         n233, n234, n235, n236, n237, n238, n239, n240, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n259, n260, n261, n262, n263,
         n264, n265, n266, n278, n286, n288, n289, n290, n291, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n311, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503;

  OAI211X1 U1 ( .A0(n376), .A1(n59), .B0(n382), .C0(n381), .Y(n383) );
  OAI21XL U2 ( .A0(n86), .A1(n39), .B0(n306), .Y(n315) );
  AOI211X1 U3 ( .A0(n311), .A1(n31), .B0(n317), .C0(n34), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n321) );
  NOR2X1 U5 ( .A(n39), .B(n83), .Y(n179) );
  OAI21XL U6 ( .A0(n2), .A1(n85), .B0(n378), .Y(n247) );
  INVXL U7 ( .A(n100), .Y(n2) );
  NOR2X1 U8 ( .A(n34), .B(n39), .Y(n289) );
  NOR2X1 U9 ( .A(n376), .B(n82), .Y(n177) );
  NAND3BX1 U10 ( .AN(n315), .B(n314), .C(n316), .Y(n320) );
  NOR2X1 U11 ( .A(n39), .B(n80), .Y(n122) );
  NAND2BX1 U12 ( .AN(n180), .B(n182), .Y(n187) );
  OAI21XL U13 ( .A0(n3), .A1(n80), .B0(n378), .Y(n141) );
  INVXL U14 ( .A(n100), .Y(n3) );
  NOR2X1 U15 ( .A(n19), .B(n101), .Y(n79) );
  NOR2X1 U16 ( .A(n17), .B(n39), .Y(n240) );
  OR2X2 U17 ( .A(n181), .B(n178), .Y(n189) );
  XOR2X2 U18 ( .A(n106), .B(n105), .Y(n374) );
  AND2X2 U19 ( .A(n80), .B(n99), .Y(n491) );
  OAI21XL U20 ( .A0(n16), .A1(n376), .B0(n378), .Y(n291) );
  NAND2BX1 U21 ( .AN(n316), .B(n317), .Y(n318) );
  NAND3X1 U22 ( .A(n181), .B(n178), .C(n180), .Y(n188) );
  XNOR2X1 U23 ( .A(n217), .B(n439), .Y(c[1]) );
  NOR2X1 U24 ( .A(n490), .B(n19), .Y(n455) );
  XOR2X2 U25 ( .A(n192), .B(n191), .Y(n259) );
  XOR2X2 U26 ( .A(n259), .B(n62), .Y(n263) );
  BUFX3 U27 ( .A(n378), .Y(n35) );
  AND2X2 U28 ( .A(n96), .B(n34), .Y(n4) );
  XNOR3X2 U29 ( .A(n235), .B(n234), .C(n233), .Y(n5) );
  XNOR3X2 U30 ( .A(n53), .B(n54), .C(n296), .Y(n6) );
  INVX1 U31 ( .A(a[12]), .Y(n39) );
  BUFX3 U32 ( .A(n59), .Y(n7) );
  INVX1 U33 ( .A(b[0]), .Y(n497) );
  BUFX3 U34 ( .A(n60), .Y(n8) );
  NAND2X1 U35 ( .A(b[0]), .B(n496), .Y(n60) );
  INVX1 U36 ( .A(n211), .Y(n9) );
  INVX1 U37 ( .A(n387), .Y(n10) );
  BUFX3 U38 ( .A(n92), .Y(n11) );
  INVX1 U39 ( .A(n388), .Y(n12) );
  INVX1 U40 ( .A(n154), .Y(n13) );
  INVX1 U41 ( .A(n222), .Y(n14) );
  INVX1 U42 ( .A(b[8]), .Y(n15) );
  INVX1 U43 ( .A(n15), .Y(n16) );
  INVX1 U44 ( .A(n15), .Y(n17) );
  INVX1 U45 ( .A(n107), .Y(n18) );
  INVX1 U46 ( .A(a[1]), .Y(n19) );
  INVX1 U47 ( .A(n19), .Y(n20) );
  INVX1 U48 ( .A(n495), .Y(n21) );
  INVX1 U49 ( .A(a[3]), .Y(n22) );
  INVXL U50 ( .A(n22), .Y(n23) );
  INVX1 U51 ( .A(a[7]), .Y(n24) );
  INVXL U52 ( .A(n24), .Y(n25) );
  INVX1 U53 ( .A(a[8]), .Y(n26) );
  INVX1 U54 ( .A(n26), .Y(n27) );
  INVX1 U55 ( .A(a[9]), .Y(n28) );
  INVX1 U56 ( .A(n28), .Y(n29) );
  INVX1 U57 ( .A(n28), .Y(n30) );
  INVX1 U58 ( .A(n101), .Y(n31) );
  OAI21XL U59 ( .A0(n102), .A1(n380), .B0(n86), .Y(n103) );
  BUFX3 U60 ( .A(b[10]), .Y(n86) );
  INVX1 U61 ( .A(n376), .Y(n32) );
  BUFX3 U62 ( .A(a[11]), .Y(n100) );
  INVX1 U63 ( .A(b[9]), .Y(n33) );
  INVX1 U64 ( .A(n33), .Y(n34) );
  XNOR3X4 U65 ( .A(n167), .B(n50), .C(n51), .Y(n260) );
  CLKINVX3 U66 ( .A(n306), .Y(n380) );
  OAI2BB1X2 U67 ( .A0N(n87), .A1N(n104), .B0(n103), .Y(n106) );
  XOR2X4 U68 ( .A(n260), .B(n168), .Y(n194) );
  OAI2BB1X1 U69 ( .A0N(n32), .A1N(n107), .B0(n35), .Y(n110) );
  OAI2BB1X1 U70 ( .A0N(n100), .A1N(n211), .B0(n35), .Y(n214) );
  AOI2BB2XL U71 ( .B0(b[0]), .B1(n380), .A0N(n35), .A1N(n377), .Y(n381) );
  OAI2BB1X1 U72 ( .A0N(n100), .A1N(n101), .B0(n378), .Y(n104) );
  NAND2BXL U73 ( .AN(a[12]), .B(n100), .Y(n378) );
  INVX1 U74 ( .A(a[10]), .Y(n36) );
  INVX1 U75 ( .A(n36), .Y(n37) );
  INVXL U76 ( .A(n36), .Y(n38) );
  AND2X1 U77 ( .A(n37), .B(n92), .Y(n105) );
  INVXL U78 ( .A(n39), .Y(n47) );
  INVX1 U79 ( .A(b[0]), .Y(n49) );
  XOR2X1 U80 ( .A(n194), .B(n169), .Y(n64) );
  XNOR3X2 U81 ( .A(n151), .B(n446), .C(n67), .Y(n50) );
  INVX1 U82 ( .A(n86), .Y(n101) );
  INVX1 U83 ( .A(n317), .Y(n314) );
  XNOR3X2 U84 ( .A(n166), .B(n165), .C(n164), .Y(n51) );
  INVXL U85 ( .A(n374), .Y(n138) );
  XNOR3X2 U86 ( .A(n52), .B(n63), .C(n216), .Y(n62) );
  XOR2X1 U87 ( .A(n210), .B(n205), .Y(n52) );
  XOR2X1 U88 ( .A(n64), .B(n447), .Y(c[2]) );
  INVXL U89 ( .A(n87), .Y(n107) );
  AOI22XL U90 ( .A0(n21), .A1(n454), .B0(n23), .B1(n453), .Y(n456) );
  AOI22XL U91 ( .A0(n27), .A1(n499), .B0(n30), .B1(n498), .Y(n501) );
  NAND2XL U92 ( .A(n85), .B(n99), .Y(n394) );
  NAND2XL U93 ( .A(n17), .B(n38), .Y(n228) );
  NAND2XL U94 ( .A(b[9]), .B(n38), .Y(n249) );
  NAND2XL U95 ( .A(n95), .B(n31), .Y(n349) );
  NAND2XL U96 ( .A(n29), .B(n92), .Y(n304) );
  NAND2XL U97 ( .A(n37), .B(n87), .Y(n303) );
  NAND2XL U98 ( .A(n92), .B(n96), .Y(n146) );
  NAND2XL U99 ( .A(a[3]), .B(n87), .Y(n145) );
  NAND2XL U100 ( .A(n97), .B(b[9]), .Y(n396) );
  NAND2XL U101 ( .A(n98), .B(n16), .Y(n397) );
  XOR2X1 U102 ( .A(n150), .B(n149), .Y(n169) );
  NAND2XL U103 ( .A(n97), .B(n86), .Y(n437) );
  NOR2X1 U104 ( .A(n226), .B(n225), .Y(n234) );
  AOI21XL U105 ( .A0(n35), .A1(n224), .B0(n387), .Y(n225) );
  NAND2XL U106 ( .A(a[7]), .B(n34), .Y(n449) );
  NAND2BXL U107 ( .AN(n84), .B(n47), .Y(n212) );
  NAND2XL U108 ( .A(n47), .B(n92), .Y(n365) );
  NAND2XL U109 ( .A(n80), .B(n38), .Y(n416) );
  NAND2XL U110 ( .A(a[7]), .B(n18), .Y(n227) );
  NAND2XL U111 ( .A(n35), .B(n305), .Y(n311) );
  NAND2BXL U112 ( .AN(b[9]), .B(n100), .Y(n305) );
  NAND2XL U113 ( .A(n31), .B(n311), .Y(n316) );
  NAND3XL U114 ( .A(n34), .B(n315), .C(n317), .Y(n319) );
  NAND2XL U115 ( .A(n95), .B(n34), .Y(n334) );
  NAND2XL U116 ( .A(n13), .B(n25), .Y(n410) );
  AOI22XL U117 ( .A0(n25), .A1(n489), .B0(n27), .B1(n488), .Y(n492) );
  NAND2XL U118 ( .A(n14), .B(n21), .Y(n66) );
  NAND2XL U119 ( .A(a[4]), .B(n9), .Y(n329) );
  NAND2XL U120 ( .A(n11), .B(a[1]), .Y(n131) );
  NAND2XL U121 ( .A(n87), .B(n96), .Y(n132) );
  NAND2XL U122 ( .A(n86), .B(a[3]), .Y(n133) );
  NAND2XL U123 ( .A(n99), .B(n31), .Y(n448) );
  NAND2XL U124 ( .A(a[3]), .B(n82), .Y(n486) );
  NAND2XL U125 ( .A(b[9]), .B(n30), .Y(n230) );
  NAND2XL U126 ( .A(n23), .B(n17), .Y(n405) );
  NAND2XL U127 ( .A(n13), .B(a[1]), .Y(n467) );
  INVXL U128 ( .A(n85), .Y(n387) );
  NAND2XL U129 ( .A(n98), .B(n92), .Y(n205) );
  NAND2XL U130 ( .A(n84), .B(n99), .Y(n413) );
  NAND2XL U131 ( .A(a[7]), .B(n86), .Y(n462) );
  NAND2XL U132 ( .A(n96), .B(n82), .Y(n477) );
  NAND2XL U133 ( .A(n29), .B(n87), .Y(n286) );
  NAND2XL U134 ( .A(n27), .B(n18), .Y(n251) );
  NAND2XL U135 ( .A(n99), .B(n92), .Y(n220) );
  NAND2XL U136 ( .A(n98), .B(n83), .Y(n350) );
  NAND2XL U137 ( .A(n95), .B(n85), .Y(n265) );
  NAND2XL U138 ( .A(n38), .B(n86), .Y(n53) );
  XNOR2X1 U139 ( .A(n288), .B(n286), .Y(n54) );
  NOR2BXL U140 ( .AN(n47), .B(n11), .Y(n108) );
  NAND2XL U141 ( .A(n12), .B(a[6]), .Y(n503) );
  NAND2XL U142 ( .A(n17), .B(n96), .Y(n347) );
  NAND2XL U143 ( .A(n97), .B(n14), .Y(n346) );
  NAND2XL U144 ( .A(n85), .B(n38), .Y(n210) );
  NAND2XL U145 ( .A(n96), .B(n12), .Y(n468) );
  NAND2XL U146 ( .A(n27), .B(n86), .Y(n221) );
  NAND2XL U147 ( .A(n99), .B(n87), .Y(n461) );
  AND2X1 U148 ( .A(n81), .B(a[1]), .Y(n202) );
  NAND2XL U149 ( .A(a[8]), .B(n92), .Y(n288) );
  INVXL U150 ( .A(n98), .Y(n385) );
  NAND2XL U151 ( .A(n85), .B(a[7]), .Y(n436) );
  NAND2XL U152 ( .A(n84), .B(n25), .Y(n395) );
  AOI22XL U153 ( .A0(n23), .A1(n458), .B0(a[4]), .B1(n457), .Y(n460) );
  XNOR3X2 U154 ( .A(n55), .B(n57), .C(n215), .Y(n216) );
  NAND2XL U155 ( .A(b[9]), .B(n27), .Y(n55) );
  NAND2XL U156 ( .A(n17), .B(n30), .Y(n57) );
  NAND2XL U157 ( .A(n34), .B(a[1]), .Y(n348) );
  NAND2XL U158 ( .A(n84), .B(n37), .Y(n173) );
  NAND2XL U159 ( .A(n16), .B(a[8]), .Y(n174) );
  NAND2XL U160 ( .A(n85), .B(n29), .Y(n175) );
  NAND2BXL U161 ( .AN(n85), .B(n47), .Y(n223) );
  NAND2BXL U162 ( .AN(n84), .B(n100), .Y(n224) );
  NAND2XL U163 ( .A(n13), .B(a[6]), .Y(n403) );
  NAND2XL U164 ( .A(n81), .B(n25), .Y(n404) );
  AOI22XL U165 ( .A0(n38), .A1(n400), .B0(n30), .B1(n399), .Y(n402) );
  NAND2XL U166 ( .A(n83), .B(a[1]), .Y(n470) );
  NAND2XL U167 ( .A(n84), .B(n95), .Y(n469) );
  NAND2XL U168 ( .A(n81), .B(n30), .Y(n418) );
  NAND2XL U169 ( .A(n82), .B(n27), .Y(n417) );
  AOI22XL U170 ( .A0(n38), .A1(n407), .B0(n32), .B1(n406), .Y(n409) );
  NAND2XL U171 ( .A(n12), .B(n27), .Y(n411) );
  XOR3X2 U172 ( .A(n58), .B(n297), .C(n359), .Y(n298) );
  NAND2XL U173 ( .A(n14), .B(n20), .Y(n58) );
  NAND2XL U174 ( .A(a[0]), .B(n11), .Y(n423) );
  INVXL U175 ( .A(n83), .Y(n211) );
  AOI22XL U176 ( .A0(a[6]), .A1(n483), .B0(n25), .B1(n482), .Y(n485) );
  NAND2XL U177 ( .A(n97), .B(n12), .Y(n487) );
  INVXL U178 ( .A(n81), .Y(n388) );
  AOI22XL U179 ( .A0(a[4]), .A1(n464), .B0(a[5]), .B1(n463), .Y(n465) );
  NAND2XL U180 ( .A(n84), .B(a[8]), .Y(n77) );
  NAND2XL U181 ( .A(n29), .B(n83), .Y(n78) );
  NAND2XL U182 ( .A(a[8]), .B(n83), .Y(n68) );
  NAND2XL U183 ( .A(n30), .B(n82), .Y(n74) );
  NAND2XL U184 ( .A(n17), .B(n20), .Y(n336) );
  NAND2XL U185 ( .A(a[3]), .B(n81), .Y(n478) );
  NAND2XL U186 ( .A(n83), .B(n25), .Y(n414) );
  XOR2X1 U187 ( .A(n254), .B(n253), .Y(n278) );
  NAND2XL U188 ( .A(n25), .B(n11), .Y(n252) );
  NAND2XL U189 ( .A(a[5]), .B(n12), .Y(n494) );
  NAND2XL U190 ( .A(n99), .B(n16), .Y(n435) );
  NAND2XL U191 ( .A(n98), .B(b[9]), .Y(n438) );
  NAND2XL U192 ( .A(n97), .B(n92), .Y(n450) );
  NAND2XL U193 ( .A(n98), .B(n87), .Y(n451) );
  NAND2XL U194 ( .A(n10), .B(n23), .Y(n351) );
  NAND2XL U195 ( .A(n95), .B(n18), .Y(n366) );
  OAI2BB1X1 U196 ( .A0N(n81), .A1N(n163), .B0(n162), .Y(n164) );
  OAI21XL U197 ( .A0(n155), .A1(n176), .B0(n82), .Y(n162) );
  AND2X1 U198 ( .A(n97), .B(n87), .Y(n67) );
  AND2X1 U199 ( .A(n37), .B(n82), .Y(n144) );
  AND2X1 U200 ( .A(n38), .B(n81), .Y(n130) );
  AND2X1 U201 ( .A(n27), .B(n80), .Y(n401) );
  AND2X1 U202 ( .A(n30), .B(n86), .Y(n250) );
  AND2X1 U203 ( .A(n95), .B(n82), .Y(n203) );
  AND2X1 U204 ( .A(n95), .B(n17), .Y(n322) );
  AND2X1 U205 ( .A(n25), .B(n80), .Y(n500) );
  INVXL U206 ( .A(n100), .Y(n376) );
  NAND2XL U207 ( .A(n10), .B(n96), .Y(n333) );
  NAND2XL U208 ( .A(n97), .B(n13), .Y(n493) );
  NAND2XL U209 ( .A(n14), .B(n23), .Y(n332) );
  NAND2XL U210 ( .A(a[6]), .B(n9), .Y(n362) );
  NAND2XL U211 ( .A(a[5]), .B(n14), .Y(n363) );
  NAND2XL U212 ( .A(a[4]), .B(n10), .Y(n364) );
  NAND2XL U213 ( .A(a[4]), .B(n17), .Y(n426) );
  NAND2XL U214 ( .A(n23), .B(n34), .Y(n425) );
  NAND2XL U215 ( .A(n13), .B(a[5]), .Y(n502) );
  NAND2XL U216 ( .A(n10), .B(n20), .Y(n300) );
  NAND2XL U217 ( .A(n23), .B(n80), .Y(n466) );
  NAND2XL U218 ( .A(n9), .B(n23), .Y(n301) );
  NAND2XL U219 ( .A(n95), .B(n9), .Y(n236) );
  NAND2XL U220 ( .A(n21), .B(n31), .Y(n428) );
  NAND2XL U221 ( .A(n20), .B(n18), .Y(n427) );
  NAND2BXL U222 ( .AN(b[1]), .B(n32), .Y(n111) );
  NAND2XL U223 ( .A(n35), .B(n111), .Y(n127) );
  INVXL U224 ( .A(b[1]), .Y(n377) );
  NAND2X1 U225 ( .A(b[1]), .B(n497), .Y(n59) );
  XNOR2X1 U226 ( .A(n138), .B(n168), .Y(n358) );
  XNOR2X1 U227 ( .A(n62), .B(n5), .Y(n302) );
  XOR2X1 U228 ( .A(n138), .B(n375), .Y(n61) );
  NAND4X1 U229 ( .A(n321), .B(n320), .C(n319), .D(n318), .Y(n384) );
  XOR2X1 U230 ( .A(n444), .B(n445), .Y(n167) );
  XOR2X1 U231 ( .A(n384), .B(n6), .Y(n361) );
  XNOR3X2 U232 ( .A(n61), .B(n169), .C(n193), .Y(n217) );
  XNOR3X2 U233 ( .A(n327), .B(n326), .C(n325), .Y(c[8]) );
  XOR2X1 U234 ( .A(n301), .B(n300), .Y(n327) );
  XOR3X2 U235 ( .A(n194), .B(n259), .C(n193), .Y(n195) );
  INVX1 U236 ( .A(n365), .Y(n375) );
  NOR2X1 U237 ( .A(n385), .B(n387), .Y(n412) );
  XNOR3X2 U238 ( .A(n219), .B(n263), .C(n217), .Y(c[4]) );
  INVX1 U239 ( .A(n368), .Y(n168) );
  XNOR3X2 U240 ( .A(n302), .B(n64), .C(n239), .Y(c[5]) );
  XOR2X1 U241 ( .A(n221), .B(n220), .Y(n235) );
  XOR3X2 U242 ( .A(n230), .B(n228), .C(n227), .Y(n233) );
  XOR2X1 U243 ( .A(n196), .B(n195), .Y(c[3]) );
  XOR3X2 U244 ( .A(n373), .B(n372), .C(n371), .Y(c[11]) );
  XOR3X2 U245 ( .A(n359), .B(n358), .C(n357), .Y(c[10]) );
  XNOR3X2 U246 ( .A(n356), .B(n355), .C(n354), .Y(n357) );
  XNOR3X2 U247 ( .A(n65), .B(n339), .C(n338), .Y(c[9]) );
  XOR2X1 U248 ( .A(n299), .B(n298), .Y(c[7]) );
  XNOR3X2 U249 ( .A(n375), .B(n260), .C(n259), .Y(n261) );
  XOR2X1 U250 ( .A(n461), .B(n462), .Y(n63) );
  XNOR3X2 U251 ( .A(n65), .B(n262), .C(n261), .Y(c[6]) );
  XOR2X1 U252 ( .A(n481), .B(n471), .Y(n262) );
  XOR2X1 U253 ( .A(n432), .B(n431), .Y(c[12]) );
  XOR2X1 U254 ( .A(n430), .B(n429), .Y(n431) );
  XOR2X1 U255 ( .A(n370), .B(n369), .Y(n371) );
  XNOR3X2 U256 ( .A(n405), .B(n4), .C(n367), .Y(n370) );
  XOR3X2 U257 ( .A(n410), .B(n368), .C(n79), .Y(n369) );
  INVX1 U258 ( .A(n181), .Y(n182) );
  INVX1 U259 ( .A(n35), .Y(n176) );
  XNOR2X1 U260 ( .A(n278), .B(n5), .Y(n65) );
  XOR2XL U261 ( .A(n278), .B(n6), .Y(n359) );
  NOR2XL U262 ( .A(n490), .B(n385), .Y(n484) );
  NOR2BX1 U263 ( .AN(a[12]), .B(n87), .Y(n102) );
  OAI21XL U264 ( .A0(n30), .A1(n377), .B0(n59), .Y(n499) );
  OAI21XL U265 ( .A0(n27), .A1(n497), .B0(n60), .Y(n498) );
  OAI21XL U266 ( .A0(n23), .A1(n377), .B0(n59), .Y(n454) );
  OAI21XL U267 ( .A0(n96), .A1(n49), .B0(n60), .Y(n453) );
  XNOR2X1 U268 ( .A(n304), .B(n303), .Y(n317) );
  AOI22X1 U269 ( .A0(n98), .A1(n473), .B0(n99), .B1(n472), .Y(n476) );
  OAI21XL U270 ( .A0(n99), .A1(n377), .B0(n59), .Y(n473) );
  OAI21XL U271 ( .A0(n98), .A1(n497), .B0(n60), .Y(n472) );
  OAI2BB1X1 U272 ( .A0N(n11), .A1N(n110), .B0(n109), .Y(n368) );
  XNOR3X2 U273 ( .A(n465), .B(n238), .C(n237), .Y(n239) );
  XOR2X1 U274 ( .A(n236), .B(n466), .Y(n237) );
  XNOR2X1 U275 ( .A(n468), .B(n467), .Y(n238) );
  OAI21XL U276 ( .A0(n30), .A1(n49), .B0(n60), .Y(n400) );
  INVXL U277 ( .A(n84), .Y(n222) );
  OAI21XL U278 ( .A0(n20), .A1(n49), .B0(n8), .Y(n440) );
  OAI21XL U279 ( .A0(n25), .A1(n49), .B0(n60), .Y(n488) );
  OAI21XL U280 ( .A0(n97), .A1(n49), .B0(n60), .Y(n463) );
  OAI21XL U281 ( .A0(n38), .A1(n49), .B0(n60), .Y(n406) );
  OAI21XL U282 ( .A0(a[6]), .A1(n49), .B0(n60), .Y(n482) );
  OAI21XL U283 ( .A0(n23), .A1(n49), .B0(n8), .Y(n457) );
  OAI21XL U284 ( .A0(n27), .A1(n496), .B0(n59), .Y(n489) );
  OAI21XL U285 ( .A0(n98), .A1(n496), .B0(n59), .Y(n464) );
  OAI21XL U286 ( .A0(n32), .A1(n377), .B0(n59), .Y(n407) );
  OAI21XL U287 ( .A0(n25), .A1(n377), .B0(n59), .Y(n483) );
  OAI21XL U288 ( .A0(n97), .A1(n377), .B0(n7), .Y(n458) );
  XNOR3X2 U289 ( .A(n437), .B(n148), .C(n147), .Y(n149) );
  XNOR3X2 U290 ( .A(n144), .B(n143), .C(n142), .Y(n150) );
  NOR2X1 U291 ( .A(n490), .B(n474), .Y(n475) );
  INVX1 U292 ( .A(n97), .Y(n474) );
  OAI21XL U293 ( .A0(n38), .A1(n377), .B0(n59), .Y(n399) );
  INVX1 U294 ( .A(n80), .Y(n490) );
  XNOR3X2 U295 ( .A(n448), .B(n449), .C(n190), .Y(n191) );
  NAND3X1 U296 ( .A(n189), .B(n188), .C(n187), .Y(n192) );
  OAI2BB1X1 U297 ( .A0N(n81), .A1N(n141), .B0(n140), .Y(n143) );
  XOR2X1 U298 ( .A(n252), .B(n251), .Y(n253) );
  XNOR3X2 U299 ( .A(n250), .B(n249), .C(n248), .Y(n254) );
  NAND2X1 U300 ( .A(n98), .B(n86), .Y(n446) );
  NOR2BX1 U301 ( .AN(n100), .B(n81), .Y(n155) );
  NAND2X1 U302 ( .A(a[7]), .B(n16), .Y(n445) );
  XOR2X1 U303 ( .A(n137), .B(n136), .Y(n193) );
  XNOR3X2 U304 ( .A(n394), .B(n135), .C(n134), .Y(n136) );
  XNOR3X2 U305 ( .A(n130), .B(n129), .C(n128), .Y(n137) );
  XNOR3X2 U306 ( .A(n374), .B(n331), .C(n330), .Y(n339) );
  XOR2X1 U307 ( .A(n329), .B(n502), .Y(n330) );
  XNOR2X1 U308 ( .A(n503), .B(n500), .Y(n331) );
  XNOR3X2 U309 ( .A(n66), .B(n492), .C(n302), .Y(n326) );
  XNOR3X2 U310 ( .A(n398), .B(n358), .C(n193), .Y(c[0]) );
  XOR2X1 U311 ( .A(n266), .B(n265), .Y(n297) );
  NAND2X1 U312 ( .A(n83), .B(n96), .Y(n266) );
  OAI2BB1X1 U313 ( .A0N(n34), .A1N(n291), .B0(n290), .Y(n296) );
  XOR2X1 U314 ( .A(n153), .B(n152), .Y(n165) );
  NAND2X1 U315 ( .A(n85), .B(a[8]), .Y(n153) );
  NAND2X1 U316 ( .A(n84), .B(n29), .Y(n152) );
  XOR2X1 U317 ( .A(n146), .B(n145), .Y(n148) );
  XOR2X1 U318 ( .A(n396), .B(n397), .Y(n135) );
  XOR3X2 U319 ( .A(n423), .B(n424), .C(n384), .Y(n432) );
  XOR2X1 U320 ( .A(n422), .B(n421), .Y(n424) );
  XOR2X1 U321 ( .A(n420), .B(n419), .Y(n421) );
  XNOR3X2 U322 ( .A(n485), .B(n264), .C(n263), .Y(n299) );
  XOR3X2 U323 ( .A(n486), .B(n487), .C(n484), .Y(n264) );
  XNOR3X2 U324 ( .A(n61), .B(n452), .C(n170), .Y(n196) );
  NOR2X1 U325 ( .A(n386), .B(n388), .Y(n452) );
  XNOR2X1 U326 ( .A(n455), .B(n456), .Y(n170) );
  XOR2X1 U327 ( .A(n418), .B(n417), .Y(n419) );
  XOR3X2 U328 ( .A(n404), .B(n403), .C(n402), .Y(n356) );
  NAND2X1 U329 ( .A(n99), .B(b[9]), .Y(n444) );
  XNOR3X2 U330 ( .A(n409), .B(n361), .C(n360), .Y(n373) );
  XNOR2X1 U331 ( .A(n408), .B(n411), .Y(n360) );
  INVX1 U332 ( .A(n82), .Y(n154) );
  NAND2BX1 U333 ( .AN(n60), .B(n47), .Y(n382) );
  XNOR3X2 U334 ( .A(n68), .B(n74), .C(n395), .Y(n128) );
  XOR3X2 U335 ( .A(n133), .B(n132), .C(n131), .Y(n134) );
  XOR2X1 U336 ( .A(n443), .B(n442), .Y(n447) );
  NOR2X1 U337 ( .A(n386), .B(n490), .Y(n442) );
  AOI22X1 U338 ( .A0(n20), .A1(n441), .B0(n21), .B1(n440), .Y(n443) );
  OAI21XL U339 ( .A0(n21), .A1(n496), .B0(n7), .Y(n441) );
  OAI2BB1X1 U340 ( .A0N(n17), .A1N(n247), .B0(n246), .Y(n248) );
  XNOR3X2 U341 ( .A(n337), .B(n336), .C(n335), .Y(n338) );
  XOR3X2 U342 ( .A(n334), .B(n333), .C(n332), .Y(n335) );
  XOR2X1 U343 ( .A(n384), .B(n501), .Y(n337) );
  AOI21X1 U344 ( .A0(n84), .A1(n214), .B0(n213), .Y(n215) );
  XOR3X2 U345 ( .A(n175), .B(n174), .C(n173), .Y(n181) );
  XOR2X1 U346 ( .A(n383), .B(n416), .Y(n420) );
  XOR2X1 U347 ( .A(n389), .B(n415), .Y(n422) );
  XOR2X1 U348 ( .A(n414), .B(n413), .Y(n415) );
  XOR3X2 U349 ( .A(n412), .B(n375), .C(n374), .Y(n389) );
  XOR2X1 U350 ( .A(n480), .B(n479), .Y(n481) );
  XOR2X1 U351 ( .A(n478), .B(n477), .Y(n479) );
  XOR2X1 U352 ( .A(n476), .B(n475), .Y(n480) );
  OAI21XL U353 ( .A0(n177), .A1(n176), .B0(n83), .Y(n178) );
  NOR2BX1 U354 ( .AN(a[12]), .B(n81), .Y(n139) );
  XOR2X1 U355 ( .A(n460), .B(n204), .Y(n219) );
  XOR3X2 U356 ( .A(n203), .B(n202), .C(n459), .Y(n204) );
  NOR2X1 U357 ( .A(n490), .B(n495), .Y(n459) );
  AND2X2 U358 ( .A(n92), .B(a[3]), .Y(n151) );
  XNOR3X2 U359 ( .A(n77), .B(n78), .C(n436), .Y(n142) );
  AND2X2 U360 ( .A(n37), .B(n83), .Y(n166) );
  XNOR2X1 U361 ( .A(n438), .B(n435), .Y(n147) );
  XNOR2X1 U362 ( .A(n450), .B(n451), .Y(n190) );
  XNOR2X1 U363 ( .A(n324), .B(n323), .Y(n325) );
  XOR2X1 U364 ( .A(n494), .B(n491), .Y(n323) );
  XNOR3X2 U365 ( .A(n322), .B(n493), .C(n361), .Y(n324) );
  XOR2X1 U366 ( .A(n353), .B(n352), .Y(n354) );
  XOR2X1 U367 ( .A(n351), .B(n350), .Y(n352) );
  XNOR3X2 U368 ( .A(n401), .B(n349), .C(n348), .Y(n353) );
  XNOR2X1 U369 ( .A(n347), .B(n346), .Y(n355) );
  NOR2BX1 U370 ( .AN(n30), .B(n490), .Y(n408) );
  NOR2X1 U371 ( .A(n386), .B(n49), .Y(n398) );
  XNOR3X2 U372 ( .A(n364), .B(n363), .C(n362), .Y(n372) );
  XOR2X1 U373 ( .A(n428), .B(n427), .Y(n429) );
  XOR2X1 U374 ( .A(n470), .B(n469), .Y(n471) );
  INVX1 U375 ( .A(n95), .Y(n386) );
  XOR2X1 U376 ( .A(n426), .B(n425), .Y(n430) );
  AOI22X1 U377 ( .A0(a[0]), .A1(n434), .B0(n20), .B1(n433), .Y(n439) );
  OAI21XL U378 ( .A0(n20), .A1(n377), .B0(n7), .Y(n434) );
  OAI21XL U379 ( .A0(n95), .A1(n49), .B0(n8), .Y(n433) );
  XOR2X1 U380 ( .A(n366), .B(n365), .Y(n367) );
  INVX1 U381 ( .A(n96), .Y(n495) );
  OAI2BB1X1 U382 ( .A0N(n80), .A1N(n127), .B0(n126), .Y(n129) );
  BUFX3 U383 ( .A(a[4]), .Y(n97) );
  BUFX3 U384 ( .A(a[6]), .Y(n99) );
  BUFX3 U385 ( .A(a[2]), .Y(n96) );
  BUFX3 U386 ( .A(a[5]), .Y(n98) );
  BUFX3 U387 ( .A(b[11]), .Y(n87) );
  BUFX3 U388 ( .A(b[3]), .Y(n81) );
  BUFX3 U389 ( .A(b[4]), .Y(n82) );
  BUFX3 U390 ( .A(b[5]), .Y(n83) );
  BUFX3 U391 ( .A(b[6]), .Y(n84) );
  BUFX3 U392 ( .A(b[7]), .Y(n85) );
  INVX1 U393 ( .A(b[1]), .Y(n496) );
  BUFX3 U394 ( .A(b[12]), .Y(n92) );
  BUFX3 U395 ( .A(a[0]), .Y(n95) );
  BUFX3 U396 ( .A(b[2]), .Y(n80) );
  OAI21XL U397 ( .A0(n108), .A1(n380), .B0(n18), .Y(n109) );
  OAI21XL U398 ( .A0(n122), .A1(n380), .B0(b[1]), .Y(n126) );
  OAI21XL U399 ( .A0(n289), .A1(n380), .B0(n17), .Y(n290) );
  OAI21XL U400 ( .A0(n179), .A1(n380), .B0(n82), .Y(n180) );
  AOI21X1 U401 ( .A0(n306), .A1(n223), .B0(n222), .Y(n226) );
  AOI21X1 U402 ( .A0(n306), .A1(n212), .B0(n211), .Y(n213) );
  OAI21XL U403 ( .A0(n240), .A1(n380), .B0(n85), .Y(n246) );
  OAI21XL U404 ( .A0(n139), .A1(n380), .B0(n80), .Y(n140) );
  OAI2BB1X1 U405 ( .A0N(a[12]), .A1N(n154), .B0(n306), .Y(n163) );
  NAND2BX4 U406 ( .AN(n100), .B(a[12]), .Y(n306) );
endmodule


module multiplier_2 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n36, n37, n38, n39, n47, n49, n50, n51, n52, n53,
         n54, n55, n57, n58, n59, n61, n63, n64, n77, n81, n83, n84, n85, n86,
         n87, n92, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n122, n127, n128, n131, n132,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n184, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n202, n203, n204, n205, n210, n211,
         n212, n213, n214, n215, n216, n217, n219, n220, n221, n225, n239,
         n240, n246, n247, n248, n249, n250, n251, n252, n253, n254, n259,
         n260, n261, n262, n263, n264, n265, n266, n286, n288, n289, n290,
         n291, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n311, n314, n315, n316, n317, n318, n319, n320, n321, n323,
         n324, n325, n326, n327, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547;

  CLKINVX3 U1 ( .A(n47), .Y(n49) );
  OAI21X1 U2 ( .A0(n388), .A1(n387), .B0(n386), .Y(n457) );
  XOR2X1 U3 ( .A(n457), .B(n458), .Y(n462) );
  OAI21XL U4 ( .A0(n107), .A1(n380), .B0(n64), .Y(n480) );
  NOR2X1 U5 ( .A(n33), .B(n99), .Y(n177) );
  NOR2X1 U6 ( .A(n8), .B(n33), .Y(n319) );
  AND2X2 U7 ( .A(n179), .B(b[3]), .Y(n385) );
  NOR2X1 U8 ( .A(n33), .B(n102), .Y(n253) );
  XNOR2X1 U9 ( .A(n288), .B(n286), .Y(n51) );
  OAI221XL U10 ( .A0(n131), .A1(n64), .B0(n63), .B1(n33), .C0(n382), .Y(n383)
         );
  NOR2XL U11 ( .A(n8), .B(n37), .Y(n334) );
  XOR3X2 U12 ( .A(n462), .B(n461), .C(n469), .Y(n472) );
  OAI21XL U13 ( .A0(n384), .A1(n180), .B0(n99), .Y(n181) );
  INVX1 U14 ( .A(n179), .Y(n384) );
  OAI21XL U15 ( .A0(b[10]), .A1(n33), .B0(n332), .Y(n336) );
  XNOR2X1 U16 ( .A(n84), .B(n500), .Y(n303) );
  XNOR3X2 U17 ( .A(n394), .B(n473), .C(n203), .Y(c[2]) );
  NAND3XL U18 ( .A(n184), .B(n178), .C(n181), .Y(n190) );
  NOR2X1 U19 ( .A(n33), .B(n98), .Y(n141) );
  XNOR3X2 U20 ( .A(n500), .B(n57), .C(n58), .Y(n498) );
  AOI21X2 U21 ( .A0(n32), .A1(n127), .B0(n122), .Y(n128) );
  CLKBUFXL U22 ( .A(n381), .Y(n1) );
  CLKBUFXL U23 ( .A(n381), .Y(n2) );
  NAND2BXL U24 ( .AN(a[12]), .B(a[11]), .Y(n381) );
  INVX1 U25 ( .A(n332), .Y(n387) );
  XOR2X1 U26 ( .A(n128), .B(n85), .Y(n149) );
  CLKINVX3 U27 ( .A(n149), .Y(n353) );
  INVX1 U28 ( .A(n246), .Y(n251) );
  NAND2BX1 U29 ( .AN(a[12]), .B(n38), .Y(n179) );
  OAI2BB1X2 U30 ( .A0N(n39), .A1N(n333), .B0(n1), .Y(n127) );
  INVX1 U31 ( .A(n37), .Y(n39) );
  INVX1 U32 ( .A(n33), .Y(n34) );
  INVX1 U33 ( .A(n38), .Y(n131) );
  INVX1 U34 ( .A(a[12]), .Y(n33) );
  XNOR3X2 U35 ( .A(n325), .B(n324), .C(n323), .Y(n3) );
  INVX1 U36 ( .A(a[11]), .Y(n37) );
  INVX1 U37 ( .A(b[3]), .Y(n4) );
  INVX1 U38 ( .A(n4), .Y(n5) );
  INVX1 U39 ( .A(b[9]), .Y(n6) );
  INVX1 U40 ( .A(n6), .Y(n7) );
  INVX1 U41 ( .A(n6), .Y(n8) );
  BUFX3 U42 ( .A(n64), .Y(n9) );
  NAND2X1 U43 ( .A(b[1]), .B(n540), .Y(n64) );
  INVX1 U44 ( .A(b[0]), .Y(n10) );
  INVX1 U45 ( .A(n211), .Y(n11) );
  INVX1 U46 ( .A(n400), .Y(n12) );
  INVX1 U47 ( .A(n397), .Y(n13) );
  BUFX3 U48 ( .A(b[4]), .Y(n14) );
  INVX1 U49 ( .A(n289), .Y(n15) );
  BUFX3 U50 ( .A(n102), .Y(n16) );
  INVX1 U51 ( .A(n538), .Y(n17) );
  INVX1 U52 ( .A(n470), .Y(n18) );
  INVX1 U53 ( .A(n506), .Y(n19) );
  INVX1 U54 ( .A(n526), .Y(n20) );
  INVX1 U55 ( .A(a[7]), .Y(n21) );
  INVXL U56 ( .A(n21), .Y(n22) );
  INVX1 U57 ( .A(a[8]), .Y(n23) );
  INVX1 U58 ( .A(n23), .Y(n24) );
  INVX1 U59 ( .A(n23), .Y(n25) );
  INVX1 U60 ( .A(a[9]), .Y(n26) );
  INVX1 U61 ( .A(n26), .Y(n27) );
  INVX1 U62 ( .A(n26), .Y(n28) );
  INVX1 U63 ( .A(a[10]), .Y(n29) );
  INVX1 U64 ( .A(n29), .Y(n30) );
  INVX1 U65 ( .A(n29), .Y(n31) );
  XOR2X1 U66 ( .A(n194), .B(n193), .Y(n246) );
  NOR2X2 U67 ( .A(n297), .B(n296), .Y(n302) );
  AOI21XL U68 ( .A0(n2), .A1(n291), .B0(n401), .Y(n296) );
  XOR2X4 U69 ( .A(n472), .B(n471), .Y(n500) );
  OAI21XL U70 ( .A0(n110), .A1(n380), .B0(n64), .Y(n505) );
  AOI22XL U71 ( .A0(n31), .A1(n410), .B0(n28), .B1(n409), .Y(n412) );
  XNOR2X1 U72 ( .A(n389), .B(n50), .Y(n57) );
  CLKINVX3 U73 ( .A(n396), .Y(n389) );
  NAND2BX1 U74 ( .AN(a[11]), .B(a[12]), .Y(n332) );
  MXI2X1 U75 ( .A(n33), .B(n385), .S0(b[4]), .Y(n388) );
  AOI21XL U76 ( .A0(n332), .A1(n290), .B0(n289), .Y(n297) );
  AOI21XL U77 ( .A0(n332), .A1(n212), .B0(n211), .Y(n213) );
  BUFX3 U78 ( .A(b[11]), .Y(n32) );
  NAND2XL U79 ( .A(a[7]), .B(b[11]), .Y(n286) );
  NOR2BXL U80 ( .AN(n34), .B(b[3]), .Y(n151) );
  NAND2BXL U81 ( .AN(n101), .B(n34), .Y(n290) );
  BUFX3 U82 ( .A(b[10]), .Y(n36) );
  INVX2 U83 ( .A(n37), .Y(n38) );
  NOR2BXL U84 ( .AN(n38), .B(b[4]), .Y(n180) );
  NAND2BXL U85 ( .AN(n100), .B(n39), .Y(n291) );
  OAI2BB1XL U86 ( .A0N(n39), .A1N(n211), .B0(n2), .Y(n214) );
  INVX1 U87 ( .A(n63), .Y(n47) );
  AOI22XL U88 ( .A0(n12), .A1(n134), .B0(n32), .B1(n132), .Y(n395) );
  NAND2X1 U89 ( .A(n24), .B(n103), .Y(n317) );
  XNOR2X1 U90 ( .A(n353), .B(n373), .Y(n378) );
  NAND2BXL U91 ( .AN(b[11]), .B(a[12]), .Y(n111) );
  NAND2BXL U92 ( .AN(n100), .B(a[12]), .Y(n212) );
  INVX1 U93 ( .A(b[10]), .Y(n333) );
  INVXL U94 ( .A(n356), .Y(n366) );
  INVX1 U95 ( .A(n247), .Y(n173) );
  XNOR2X1 U96 ( .A(n315), .B(n50), .Y(n84) );
  XOR2X1 U97 ( .A(n315), .B(n3), .Y(n356) );
  NAND2XL U98 ( .A(n187), .B(n182), .Y(n191) );
  AOI21X1 U99 ( .A0(n332), .A1(n111), .B0(n333), .Y(n122) );
  NAND2X1 U100 ( .A(n101), .B(n27), .Y(n176) );
  NAND2X1 U101 ( .A(n102), .B(n24), .Y(n175) );
  AOI21X1 U102 ( .A0(n100), .A1(n214), .B0(n213), .Y(n240) );
  NAND2XL U103 ( .A(n107), .B(n5), .Y(n510) );
  NAND2XL U104 ( .A(n108), .B(n5), .Y(n519) );
  AOI22X1 U105 ( .A0(n22), .A1(n525), .B0(n25), .B1(n524), .Y(n529) );
  INVXL U106 ( .A(n378), .Y(n202) );
  XOR3X2 U107 ( .A(n51), .B(n302), .C(n301), .Y(n50) );
  NOR2XL U108 ( .A(n397), .B(n401), .Y(n424) );
  XOR2X1 U109 ( .A(n402), .B(n523), .Y(n535) );
  NAND2X1 U110 ( .A(n188), .B(n187), .Y(n189) );
  NOR2XL U111 ( .A(n398), .B(n401), .Y(n520) );
  XOR3X2 U112 ( .A(n52), .B(n411), .C(n53), .Y(n365) );
  XOR3X2 U113 ( .A(n412), .B(n358), .C(n357), .Y(n52) );
  XNOR3X2 U114 ( .A(n364), .B(n363), .C(n362), .Y(n53) );
  XOR2X1 U115 ( .A(n173), .B(n452), .Y(c[1]) );
  XOR3X2 U116 ( .A(n377), .B(n54), .C(n376), .Y(c[11]) );
  XOR3X2 U117 ( .A(n372), .B(n371), .C(n370), .Y(n54) );
  XOR3X2 U118 ( .A(n355), .B(n84), .C(n55), .Y(c[9]) );
  XNOR3X2 U119 ( .A(n354), .B(n353), .C(n352), .Y(n55) );
  NOR2XL U120 ( .A(n399), .B(n4), .Y(n478) );
  NAND2XL U121 ( .A(n101), .B(n110), .Y(n404) );
  NAND2XL U122 ( .A(n7), .B(n31), .Y(n261) );
  NAND2XL U123 ( .A(b[7]), .B(n107), .Y(n358) );
  NAND2XL U124 ( .A(n16), .B(n17), .Y(n363) );
  NAND2XL U125 ( .A(n101), .B(n25), .Y(n459) );
  AOI22XL U126 ( .A0(n25), .A1(n542), .B0(n28), .B1(n541), .Y(n544) );
  NAND2XL U127 ( .A(n108), .B(n7), .Y(n406) );
  NAND2XL U128 ( .A(n109), .B(n102), .Y(n407) );
  NAND2XL U129 ( .A(n11), .B(n106), .Y(n314) );
  NAND2XL U130 ( .A(n104), .B(b[7]), .Y(n311) );
  OAI21XL U131 ( .A0(n334), .A1(n384), .B0(n36), .Y(n335) );
  INVXL U132 ( .A(n101), .Y(n401) );
  NAND2XL U133 ( .A(n22), .B(n12), .Y(n264) );
  NAND2XL U134 ( .A(n34), .B(n12), .Y(n249) );
  NAND2XL U135 ( .A(n2), .B(n318), .Y(n321) );
  NAND2BXL U136 ( .AN(n102), .B(n39), .Y(n318) );
  NAND2XL U137 ( .A(a[7]), .B(n8), .Y(n475) );
  OAI2BB1X1 U138 ( .A0N(n5), .A1N(n153), .B0(n152), .Y(n163) );
  NAND2XL U139 ( .A(n2), .B(n150), .Y(n153) );
  NAND2BXL U140 ( .AN(n98), .B(n38), .Y(n150) );
  NAND2XL U141 ( .A(n14), .B(n22), .Y(n422) );
  NAND2XL U142 ( .A(n19), .B(b[7]), .Y(n372) );
  NAND2XL U143 ( .A(n98), .B(n31), .Y(n428) );
  NAND2XL U144 ( .A(n31), .B(b[3]), .Y(n146) );
  NAND2XL U145 ( .A(n107), .B(n14), .Y(n518) );
  NAND2XL U146 ( .A(n110), .B(n36), .Y(n474) );
  NAND2XL U147 ( .A(n18), .B(n16), .Y(n416) );
  NAND2XL U148 ( .A(n100), .B(n20), .Y(n425) );
  NAND2XL U149 ( .A(n101), .B(n106), .Y(n349) );
  NAND2XL U150 ( .A(n14), .B(n25), .Y(n429) );
  NAND2XL U151 ( .A(n110), .B(n7), .Y(n463) );
  NAND2XL U152 ( .A(n16), .B(n105), .Y(n338) );
  NAND2XL U153 ( .A(n110), .B(b[11]), .Y(n487) );
  NAND2XL U154 ( .A(n15), .B(n104), .Y(n501) );
  NAND2XL U155 ( .A(n108), .B(n14), .Y(n530) );
  NAND2XL U156 ( .A(n27), .B(b[11]), .Y(n316) );
  NAND2XL U157 ( .A(n108), .B(b[11]), .Y(n465) );
  NAND2XL U158 ( .A(n25), .B(n32), .Y(n263) );
  XOR2X1 U159 ( .A(n221), .B(n220), .Y(n225) );
  NAND2XL U160 ( .A(n30), .B(n103), .Y(n85) );
  NAND2XL U161 ( .A(n99), .B(n30), .Y(n458) );
  NAND2XL U162 ( .A(n103), .B(n106), .Y(n166) );
  NAND2XL U163 ( .A(n107), .B(n32), .Y(n165) );
  NAND2XL U164 ( .A(n17), .B(n8), .Y(n415) );
  NAND2XL U165 ( .A(n104), .B(n8), .Y(n350) );
  NAND2XL U166 ( .A(n99), .B(n105), .Y(n502) );
  NAND2XL U167 ( .A(a[7]), .B(b[10]), .Y(n488) );
  NAND2XL U168 ( .A(n2), .B(n252), .Y(n259) );
  NAND2XL U169 ( .A(n108), .B(n15), .Y(n359) );
  NAND2XL U170 ( .A(n8), .B(n105), .Y(n361) );
  NAND2XL U171 ( .A(n101), .B(n22), .Y(n449) );
  NAND2XL U172 ( .A(n100), .B(a[7]), .Y(n405) );
  NAND2XL U173 ( .A(n5), .B(n22), .Y(n414) );
  NAND2XL U174 ( .A(n14), .B(n20), .Y(n413) );
  NAND2XL U175 ( .A(n13), .B(n11), .Y(n357) );
  NAND2XL U176 ( .A(n100), .B(n31), .Y(n174) );
  NAND2XL U177 ( .A(n5), .B(n110), .Y(n546) );
  NAND2XL U178 ( .A(n14), .B(n109), .Y(n545) );
  NAND2XL U179 ( .A(n5), .B(n28), .Y(n430) );
  NAND2XL U180 ( .A(a[7]), .B(n102), .Y(n464) );
  NAND2XL U181 ( .A(n106), .B(n14), .Y(n509) );
  NAND2XL U182 ( .A(n101), .B(n30), .Y(n216) );
  NAND2XL U183 ( .A(n102), .B(n28), .Y(n215) );
  AOI22XL U184 ( .A0(n31), .A1(n419), .B0(n39), .B1(n418), .Y(n421) );
  NAND2XL U185 ( .A(n5), .B(n25), .Y(n423) );
  NAND2XL U186 ( .A(n100), .B(n107), .Y(n339) );
  XNOR3X2 U187 ( .A(n395), .B(n497), .C(n394), .Y(n58) );
  XOR3X2 U188 ( .A(n86), .B(n87), .C(n59), .Y(n210) );
  NOR2X1 U189 ( .A(n527), .B(n538), .Y(n59) );
  AOI22XL U190 ( .A0(n20), .A1(n515), .B0(n22), .B1(n514), .Y(n517) );
  NAND2XL U191 ( .A(n100), .B(n24), .Y(n92) );
  NAND2XL U192 ( .A(n28), .B(n99), .Y(n95) );
  NAND2XL U193 ( .A(n103), .B(n105), .Y(n135) );
  NAND2XL U194 ( .A(n32), .B(n106), .Y(n136) );
  NAND2XL U195 ( .A(n24), .B(n99), .Y(n96) );
  NAND2XL U196 ( .A(n27), .B(b[4]), .Y(n97) );
  INVXL U197 ( .A(n110), .Y(n526) );
  NAND2XL U198 ( .A(n99), .B(n22), .Y(n426) );
  XNOR2XL U199 ( .A(n435), .B(n547), .Y(n436) );
  NAND2XL U200 ( .A(n104), .B(n12), .Y(n435) );
  NAND2XL U201 ( .A(n32), .B(n31), .Y(n417) );
  NAND2XL U202 ( .A(n108), .B(n103), .Y(n476) );
  NAND2XL U203 ( .A(n109), .B(n32), .Y(n477) );
  NAND2XL U204 ( .A(n109), .B(n8), .Y(n451) );
  NAND2XL U205 ( .A(n110), .B(n102), .Y(n448) );
  INVXL U206 ( .A(n100), .Y(n289) );
  INVXL U207 ( .A(n103), .Y(n400) );
  AND2X1 U208 ( .A(n31), .B(b[4]), .Y(n164) );
  XNOR3X2 U209 ( .A(n61), .B(n417), .C(n337), .Y(n547) );
  NAND2XL U210 ( .A(n28), .B(n103), .Y(n61) );
  AND2X1 U211 ( .A(n15), .B(n105), .Y(n327) );
  AND2X1 U212 ( .A(n27), .B(n36), .Y(n262) );
  AND2X1 U213 ( .A(n108), .B(n99), .Y(n346) );
  INVX1 U214 ( .A(n178), .Y(n182) );
  OAI21XL U215 ( .A0(n177), .A1(n387), .B0(n14), .Y(n178) );
  AND2X1 U216 ( .A(n30), .B(b[10]), .Y(n325) );
  AND2X1 U217 ( .A(n22), .B(n98), .Y(n543) );
  INVX1 U218 ( .A(n181), .Y(n188) );
  XOR2X1 U219 ( .A(n460), .B(n459), .Y(n461) );
  NAND2XL U220 ( .A(n100), .B(n28), .Y(n460) );
  NAND2XL U221 ( .A(n109), .B(n103), .Y(n219) );
  NAND2XL U222 ( .A(n7), .B(n24), .Y(n217) );
  NAND2XL U223 ( .A(n107), .B(n99), .Y(n522) );
  NAND2XL U224 ( .A(n15), .B(n106), .Y(n521) );
  NAND2XL U225 ( .A(n13), .B(n15), .Y(n371) );
  NAND2XL U226 ( .A(n104), .B(n32), .Y(n375) );
  NAND2XL U227 ( .A(n18), .B(n8), .Y(n438) );
  NAND2XL U228 ( .A(n14), .B(n105), .Y(n493) );
  NAND2XL U229 ( .A(a[1]), .B(n32), .Y(n440) );
  AND2X1 U230 ( .A(n25), .B(n98), .Y(n411) );
  AND2X1 U231 ( .A(n16), .B(a[0]), .Y(n536) );
  NAND2XL U232 ( .A(n20), .B(n11), .Y(n370) );
  NAND2XL U233 ( .A(n19), .B(n16), .Y(n439) );
  NAND2XL U234 ( .A(b[0]), .B(n539), .Y(n63) );
  NAND2XL U235 ( .A(n2), .B(n140), .Y(n143) );
  NAND2BXL U236 ( .AN(b[1]), .B(n39), .Y(n140) );
  AOI2BB2XL U237 ( .B0(b[0]), .B1(n387), .A0N(n2), .A1N(n380), .Y(n382) );
  INVXL U238 ( .A(b[1]), .Y(n380) );
  XOR2X1 U239 ( .A(n149), .B(n395), .Y(n367) );
  XOR2X1 U240 ( .A(n547), .B(n3), .Y(n369) );
  XOR2X1 U241 ( .A(n246), .B(n389), .Y(n305) );
  XNOR3X2 U242 ( .A(n202), .B(n195), .C(n394), .Y(n247) );
  XOR3X2 U243 ( .A(n300), .B(n299), .C(n298), .Y(n301) );
  XOR3X2 U244 ( .A(n369), .B(n536), .C(n537), .Y(c[8]) );
  XNOR3X2 U245 ( .A(n202), .B(n251), .C(n195), .Y(n204) );
  XNOR2X1 U246 ( .A(n500), .B(n395), .Y(n203) );
  XOR3X2 U247 ( .A(n520), .B(n50), .C(n396), .Y(n402) );
  XNOR3X2 U248 ( .A(n251), .B(n513), .C(n250), .Y(n304) );
  XOR2X1 U249 ( .A(n249), .B(n503), .Y(n250) );
  XOR2X1 U250 ( .A(n512), .B(n511), .Y(n513) );
  XOR2X1 U251 ( .A(n502), .B(n501), .Y(n503) );
  XNOR3X2 U252 ( .A(n305), .B(n248), .C(n247), .Y(c[4]) );
  XOR2X1 U253 ( .A(n486), .B(n210), .Y(n248) );
  XOR2X1 U254 ( .A(n499), .B(n498), .Y(c[5]) );
  XNOR3X2 U255 ( .A(n77), .B(n81), .C(n83), .Y(n376) );
  XNOR2XL U256 ( .A(n395), .B(n373), .Y(n77) );
  XNOR2X1 U257 ( .A(n415), .B(n416), .Y(n81) );
  XOR3X2 U258 ( .A(n422), .B(n375), .C(n374), .Y(n83) );
  INVX1 U259 ( .A(n249), .Y(n373) );
  XNOR3X2 U260 ( .A(n205), .B(n204), .C(n203), .Y(c[3]) );
  XOR2X1 U261 ( .A(n483), .B(n478), .Y(n205) );
  XNOR3X2 U262 ( .A(n367), .B(n366), .C(n365), .Y(c[10]) );
  XOR2X1 U263 ( .A(n331), .B(n330), .Y(c[7]) );
  XNOR3X2 U264 ( .A(n327), .B(n326), .C(n356), .Y(n330) );
  XOR2X1 U265 ( .A(n304), .B(n303), .Y(c[6]) );
  XOR2X1 U266 ( .A(n445), .B(n444), .Y(c[12]) );
  XOR2X1 U267 ( .A(n535), .B(n534), .Y(n537) );
  XOR2X1 U268 ( .A(n533), .B(n532), .Y(n534) );
  XOR2X1 U269 ( .A(n531), .B(n530), .Y(n532) );
  INVX1 U270 ( .A(n184), .Y(n187) );
  NOR2X1 U271 ( .A(n527), .B(n397), .Y(n516) );
  OAI21XL U272 ( .A0(n32), .A1(n131), .B0(n2), .Y(n134) );
  OAI2BB1X1 U273 ( .A0N(n38), .A1N(b[4]), .B0(n4), .Y(n386) );
  AOI22X1 U274 ( .A0(n18), .A1(n485), .B0(n19), .B1(n484), .Y(n486) );
  OAI21XL U275 ( .A0(n19), .A1(n380), .B0(n9), .Y(n485) );
  OAI21XL U276 ( .A0(n18), .A1(n540), .B0(n49), .Y(n484) );
  OAI21XL U277 ( .A0(n31), .A1(n380), .B0(n64), .Y(n409) );
  OAI21XL U278 ( .A0(n28), .A1(n10), .B0(n49), .Y(n410) );
  OAI2BB1X1 U279 ( .A0N(n8), .A1N(n336), .B0(n335), .Y(n337) );
  OAI21XL U280 ( .A0(n25), .A1(n380), .B0(n64), .Y(n525) );
  OAI21XL U281 ( .A0(n39), .A1(n380), .B0(n64), .Y(n419) );
  OAI21XL U282 ( .A0(n22), .A1(n380), .B0(n64), .Y(n515) );
  OAI21XL U283 ( .A0(n109), .A1(n10), .B0(n63), .Y(n504) );
  OAI21XL U284 ( .A0(n22), .A1(n10), .B0(n49), .Y(n524) );
  OAI21XL U285 ( .A0(n106), .A1(n10), .B0(n49), .Y(n479) );
  OAI21XL U286 ( .A0(n105), .A1(n540), .B0(n49), .Y(n453) );
  OAI21XL U287 ( .A0(n31), .A1(n10), .B0(n49), .Y(n418) );
  OAI21XL U288 ( .A0(n20), .A1(n10), .B0(n49), .Y(n514) );
  AOI22X1 U289 ( .A0(n19), .A1(n490), .B0(n13), .B1(n489), .Y(n491) );
  OAI21XL U290 ( .A0(n13), .A1(n380), .B0(n64), .Y(n490) );
  OAI21XL U291 ( .A0(n108), .A1(n10), .B0(n49), .Y(n489) );
  INVX1 U292 ( .A(n98), .Y(n527) );
  XOR2X1 U293 ( .A(n170), .B(n169), .Y(n394) );
  XNOR3X2 U294 ( .A(n450), .B(n168), .C(n167), .Y(n169) );
  XNOR3X2 U295 ( .A(n164), .B(n163), .C(n162), .Y(n170) );
  NAND2X1 U296 ( .A(n108), .B(n36), .Y(n450) );
  XOR2X1 U297 ( .A(n148), .B(n147), .Y(n195) );
  XNOR3X2 U298 ( .A(n404), .B(n139), .C(n138), .Y(n148) );
  XNOR3X2 U299 ( .A(n146), .B(n145), .C(n144), .Y(n147) );
  XOR3X2 U300 ( .A(n176), .B(n175), .C(n174), .Y(n184) );
  XNOR3X2 U301 ( .A(n240), .B(n239), .C(n225), .Y(n396) );
  XNOR2X1 U302 ( .A(n488), .B(n487), .Y(n239) );
  XNOR3X2 U303 ( .A(n474), .B(n475), .C(n192), .Y(n193) );
  NAND3X1 U304 ( .A(n191), .B(n190), .C(n189), .Y(n194) );
  XOR2X1 U305 ( .A(n266), .B(n265), .Y(n315) );
  XOR2X1 U306 ( .A(n264), .B(n263), .Y(n265) );
  XNOR3X2 U307 ( .A(n262), .B(n261), .C(n260), .Y(n266) );
  NOR2X1 U308 ( .A(n400), .B(n470), .Y(n471) );
  INVX1 U309 ( .A(n107), .Y(n470) );
  NAND2X1 U310 ( .A(n110), .B(n103), .Y(n299) );
  OAI21XL U311 ( .A0(n151), .A1(n387), .B0(n98), .Y(n152) );
  XNOR2X1 U312 ( .A(n216), .B(n215), .Y(n221) );
  XOR2X1 U313 ( .A(n510), .B(n509), .Y(n511) );
  NOR2BX1 U314 ( .AN(n28), .B(n527), .Y(n420) );
  NAND2X1 U315 ( .A(n104), .B(n14), .Y(n86) );
  NAND2X1 U316 ( .A(n5), .B(n105), .Y(n87) );
  AND2X2 U317 ( .A(n11), .B(n104), .Y(n497) );
  XNOR3X2 U318 ( .A(n408), .B(n367), .C(n195), .Y(c[0]) );
  NOR2X1 U319 ( .A(n399), .B(n10), .Y(n408) );
  XOR2X1 U320 ( .A(n456), .B(n455), .Y(n473) );
  NOR2X1 U321 ( .A(n399), .B(n527), .Y(n455) );
  AOI22X1 U322 ( .A0(n105), .A1(n454), .B0(n17), .B1(n453), .Y(n456) );
  OAI21XL U323 ( .A0(n106), .A1(n380), .B0(n9), .Y(n454) );
  XOR2X1 U324 ( .A(n166), .B(n165), .Y(n168) );
  XOR2X1 U325 ( .A(n406), .B(n407), .Y(n139) );
  XNOR3X2 U326 ( .A(n517), .B(n306), .C(n305), .Y(n331) );
  XOR3X2 U327 ( .A(n518), .B(n519), .C(n516), .Y(n306) );
  XOR2X1 U328 ( .A(n219), .B(n217), .Y(n220) );
  XOR2X1 U329 ( .A(n468), .B(n467), .Y(n469) );
  XOR2X1 U330 ( .A(n464), .B(n463), .Y(n468) );
  XOR2X1 U331 ( .A(n466), .B(n465), .Y(n467) );
  XOR2X1 U332 ( .A(n432), .B(n431), .Y(n433) );
  XOR2X1 U333 ( .A(n430), .B(n429), .Y(n431) );
  XOR2X1 U334 ( .A(n383), .B(n428), .Y(n432) );
  XOR3X2 U335 ( .A(n545), .B(n546), .C(n351), .Y(n354) );
  XOR2X1 U336 ( .A(n350), .B(n349), .Y(n351) );
  NAND2X1 U337 ( .A(n102), .B(n30), .Y(n288) );
  XNOR3X2 U338 ( .A(n421), .B(n369), .C(n368), .Y(n377) );
  XNOR2X1 U339 ( .A(n420), .B(n423), .Y(n368) );
  NAND2X1 U340 ( .A(n109), .B(n36), .Y(n466) );
  XNOR3X2 U341 ( .A(n348), .B(n347), .C(n547), .Y(n355) );
  XOR2X1 U342 ( .A(n339), .B(n338), .Y(n348) );
  XOR2X1 U343 ( .A(n543), .B(n346), .Y(n347) );
  NAND2X1 U344 ( .A(n25), .B(n36), .Y(n298) );
  OAI2BB1X1 U345 ( .A0N(n8), .A1N(n321), .B0(n320), .Y(n323) );
  OAI21XL U346 ( .A0(n319), .A1(n387), .B0(n16), .Y(n320) );
  XNOR3X2 U347 ( .A(n92), .B(n95), .C(n449), .Y(n162) );
  XNOR3X2 U348 ( .A(n96), .B(n97), .C(n405), .Y(n144) );
  XOR3X2 U349 ( .A(n361), .B(n360), .C(n359), .Y(n362) );
  NAND2X1 U350 ( .A(n104), .B(n36), .Y(n360) );
  XOR2X1 U351 ( .A(n317), .B(n316), .Y(n324) );
  XNOR3X2 U352 ( .A(n137), .B(n136), .C(n135), .Y(n138) );
  NAND2X1 U353 ( .A(n36), .B(n107), .Y(n137) );
  NAND2X1 U354 ( .A(n7), .B(n27), .Y(n300) );
  OAI2BB1X1 U355 ( .A0N(n102), .A1N(n259), .B0(n254), .Y(n260) );
  OAI21XL U356 ( .A0(n253), .A1(n387), .B0(n101), .Y(n254) );
  NAND2BXL U357 ( .AN(n101), .B(n39), .Y(n252) );
  XOR2X1 U358 ( .A(n508), .B(n507), .Y(n512) );
  NOR2X1 U359 ( .A(n527), .B(n506), .Y(n507) );
  AOI22X1 U360 ( .A0(n109), .A1(n505), .B0(n110), .B1(n504), .Y(n508) );
  INVX1 U361 ( .A(n108), .Y(n506) );
  XOR2X1 U362 ( .A(n529), .B(n528), .Y(n533) );
  NOR2X1 U363 ( .A(n527), .B(n526), .Y(n528) );
  XOR2X1 U364 ( .A(n482), .B(n481), .Y(n483) );
  NOR2X1 U365 ( .A(n398), .B(n527), .Y(n481) );
  AOI22X1 U366 ( .A0(n106), .A1(n480), .B0(n107), .B1(n479), .Y(n482) );
  XOR2X1 U367 ( .A(n437), .B(n436), .Y(n445) );
  XOR2X1 U368 ( .A(n434), .B(n433), .Y(n437) );
  XOR2X1 U369 ( .A(n403), .B(n427), .Y(n434) );
  XOR2X1 U370 ( .A(n426), .B(n425), .Y(n427) );
  XOR2X1 U371 ( .A(n378), .B(n424), .Y(n403) );
  XOR2X1 U372 ( .A(n496), .B(n495), .Y(n499) );
  XOR2X1 U373 ( .A(n494), .B(n493), .Y(n495) );
  XOR2X1 U374 ( .A(n492), .B(n491), .Y(n496) );
  NAND2X1 U375 ( .A(n17), .B(n5), .Y(n494) );
  XOR2X1 U376 ( .A(n414), .B(n413), .Y(n364) );
  INVX1 U377 ( .A(n105), .Y(n398) );
  INVX1 U378 ( .A(n109), .Y(n397) );
  XNOR2X1 U379 ( .A(n476), .B(n477), .Y(n192) );
  XNOR2X1 U380 ( .A(n451), .B(n448), .Y(n167) );
  INVX1 U381 ( .A(n544), .Y(n352) );
  OAI21XL U382 ( .A0(n28), .A1(n539), .B0(n9), .Y(n542) );
  OAI21XL U383 ( .A0(n25), .A1(n10), .B0(n49), .Y(n541) );
  INVX1 U384 ( .A(n99), .Y(n211) );
  AOI22X1 U385 ( .A0(a[0]), .A1(n447), .B0(a[1]), .B1(n446), .Y(n452) );
  OAI21XL U386 ( .A0(a[1]), .A1(n539), .B0(n9), .Y(n447) );
  OAI21XL U387 ( .A0(n104), .A1(n10), .B0(n49), .Y(n446) );
  XOR2X1 U388 ( .A(n314), .B(n311), .Y(n326) );
  XOR2X1 U389 ( .A(n522), .B(n521), .Y(n523) );
  XOR2X1 U390 ( .A(n443), .B(n442), .Y(n444) );
  XOR2X1 U391 ( .A(n439), .B(n438), .Y(n443) );
  XOR2X1 U392 ( .A(n441), .B(n440), .Y(n442) );
  NAND2X1 U393 ( .A(n109), .B(n5), .Y(n531) );
  NAND2X1 U394 ( .A(n17), .B(n36), .Y(n441) );
  NAND2X1 U395 ( .A(n18), .B(n98), .Y(n492) );
  INVX1 U396 ( .A(n104), .Y(n399) );
  NAND2X1 U397 ( .A(a[1]), .B(n36), .Y(n374) );
  INVX1 U398 ( .A(n106), .Y(n538) );
  OAI2BB1X1 U399 ( .A0N(n98), .A1N(n143), .B0(n142), .Y(n145) );
  OAI21XL U400 ( .A0(n141), .A1(n387), .B0(b[1]), .Y(n142) );
  BUFX3 U401 ( .A(a[3]), .Y(n107) );
  BUFX3 U402 ( .A(a[6]), .Y(n110) );
  BUFX3 U403 ( .A(a[2]), .Y(n106) );
  BUFX3 U404 ( .A(a[4]), .Y(n108) );
  BUFX3 U405 ( .A(a[5]), .Y(n109) );
  BUFX3 U406 ( .A(b[6]), .Y(n100) );
  BUFX3 U407 ( .A(b[8]), .Y(n102) );
  BUFX3 U408 ( .A(a[1]), .Y(n105) );
  INVX1 U409 ( .A(b[0]), .Y(n540) );
  BUFX3 U410 ( .A(b[12]), .Y(n103) );
  BUFX3 U411 ( .A(b[7]), .Y(n101) );
  BUFX3 U412 ( .A(b[5]), .Y(n99) );
  INVX1 U413 ( .A(b[1]), .Y(n539) );
  BUFX3 U414 ( .A(b[2]), .Y(n98) );
  BUFX3 U415 ( .A(a[0]), .Y(n104) );
  OAI21XL U416 ( .A0(n103), .A1(n33), .B0(n332), .Y(n132) );
endmodule


module multiplier_1 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n43, n47, n49, n50,
         n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n72, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n92, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n122, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n202, n203, n204, n205, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n230, n233, n234, n235, n236, n237, n238, n239, n240,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n259, n260,
         n261, n262, n263, n264, n265, n266, n278, n286, n288, n289, n290,
         n291, n292, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n343, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489;

  CLKINVX3 U1 ( .A(n16), .Y(n17) );
  XOR2X1 U2 ( .A(n177), .B(n176), .Y(n187) );
  INVX1 U3 ( .A(n262), .Y(n216) );
  OAI221XL U4 ( .A0(n1), .A1(n55), .B0(n373), .B1(n54), .C0(n376), .Y(n377) );
  INVX1 U5 ( .A(n36), .Y(n1) );
  NAND2X1 U6 ( .A(n86), .B(n101), .Y(n176) );
  NOR2BX1 U7 ( .AN(n96), .B(n480), .Y(n444) );
  NOR2X1 U8 ( .A(n32), .B(n10), .Y(n107) );
  NAND2XL U9 ( .A(n17), .B(n99), .Y(n387) );
  XNOR3X2 U10 ( .A(n359), .B(n263), .C(n262), .Y(n264) );
  OAI2BB1XL U11 ( .A0N(n16), .A1N(n37), .B0(n374), .Y(n290) );
  XOR2X1 U12 ( .A(n62), .B(n429), .Y(c[1]) );
  NAND2BX1 U13 ( .AN(n103), .B(n102), .Y(n374) );
  OAI21X1 U14 ( .A0(n104), .A1(n375), .B0(n87), .Y(n105) );
  INVX2 U15 ( .A(n371), .Y(n140) );
  AND2X2 U16 ( .A(n85), .B(n33), .Y(n188) );
  OAI2BB1X1 U17 ( .A0N(n36), .A1N(n303), .B0(n302), .Y(n314) );
  CLKINVX3 U18 ( .A(n302), .Y(n375) );
  NAND2BX2 U19 ( .AN(n102), .B(n103), .Y(n302) );
  BUFX4 U20 ( .A(a[11]), .Y(n102) );
  XOR2X1 U21 ( .A(n190), .B(n189), .Y(n262) );
  XNOR3X2 U22 ( .A(n237), .B(n236), .C(n235), .Y(n2) );
  XNOR3X2 U23 ( .A(n40), .B(n43), .C(n291), .Y(n3) );
  XNOR2X1 U24 ( .A(n433), .B(n432), .Y(n4) );
  NAND2XL U25 ( .A(b[0]), .B(n484), .Y(n5) );
  INVX1 U26 ( .A(n178), .Y(n6) );
  INVX1 U27 ( .A(n210), .Y(n7) );
  INVX1 U28 ( .A(n382), .Y(n8) );
  INVX1 U29 ( .A(n303), .Y(n9) );
  INVX1 U30 ( .A(b[12]), .Y(n10) );
  INVX1 U31 ( .A(n10), .Y(n11) );
  INVX1 U32 ( .A(n10), .Y(n12) );
  INVX1 U33 ( .A(n380), .Y(n13) );
  INVX1 U34 ( .A(n99), .Y(n380) );
  INVX1 U35 ( .A(b[0]), .Y(n14) );
  INVX1 U36 ( .A(n224), .Y(n15) );
  INVX1 U37 ( .A(b[8]), .Y(n16) );
  INVXL U38 ( .A(n16), .Y(n18) );
  INVX1 U39 ( .A(b[9]), .Y(n19) );
  INVX1 U40 ( .A(n19), .Y(n20) );
  INVX1 U41 ( .A(n109), .Y(n21) );
  INVX1 U42 ( .A(n483), .Y(n22) );
  INVX1 U43 ( .A(a[3]), .Y(n23) );
  INVXL U44 ( .A(n23), .Y(n24) );
  INVX1 U45 ( .A(n463), .Y(n25) );
  INVX1 U46 ( .A(n479), .Y(n26) );
  INVX1 U47 ( .A(a[7]), .Y(n27) );
  INVX1 U48 ( .A(n27), .Y(n28) );
  INVX1 U49 ( .A(a[8]), .Y(n29) );
  INVX1 U50 ( .A(n29), .Y(n30) );
  INVX1 U51 ( .A(n398), .Y(n31) );
  INVX1 U52 ( .A(a[10]), .Y(n32) );
  INVX1 U53 ( .A(n32), .Y(n33) );
  INVX1 U54 ( .A(n32), .Y(n34) );
  NAND2X1 U55 ( .A(a[8]), .B(n84), .Y(n67) );
  NAND2X1 U56 ( .A(n87), .B(a[3]), .Y(n135) );
  XOR2X2 U57 ( .A(n153), .B(n152), .Y(n174) );
  CLKINVX3 U58 ( .A(n263), .Y(n193) );
  NAND2XL U59 ( .A(n6), .B(n13), .Y(n489) );
  AOI22XL U60 ( .A0(n25), .A1(n453), .B0(n13), .B1(n452), .Y(n454) );
  NAND2XL U61 ( .A(n13), .B(n84), .Y(n348) );
  AND2X1 U62 ( .A(n99), .B(n82), .Y(n65) );
  AOI22XL U63 ( .A0(n99), .A1(n462), .B0(n100), .B1(n461), .Y(n465) );
  NAND2XL U64 ( .A(n99), .B(b[9]), .Y(n428) );
  BUFX3 U65 ( .A(n374), .Y(n81) );
  INVX1 U66 ( .A(b[1]), .Y(n35) );
  BUFX3 U67 ( .A(n103), .Y(n36) );
  BUFX3 U68 ( .A(a[11]), .Y(n37) );
  NAND2XL U69 ( .A(b[1]), .B(n485), .Y(n38) );
  NAND2XL U70 ( .A(n85), .B(n101), .Y(n155) );
  NAND2XL U71 ( .A(b[1]), .B(n485), .Y(n54) );
  NAND2XL U72 ( .A(n86), .B(a[8]), .Y(n162) );
  OAI2BB1XL U73 ( .A0N(n37), .A1N(n109), .B0(n81), .Y(n122) );
  OAI2BB1XL U74 ( .A0N(n37), .A1N(n178), .B0(n81), .Y(n181) );
  BUFX3 U75 ( .A(a[5]), .Y(n99) );
  BUFX3 U76 ( .A(a[2]), .Y(n97) );
  BUFX3 U77 ( .A(a[12]), .Y(n103) );
  NAND2XL U78 ( .A(n81), .B(n141), .Y(n144) );
  NAND2XL U79 ( .A(n97), .B(b[3]), .Y(n457) );
  NAND2XL U80 ( .A(n85), .B(n97), .Y(n318) );
  NAND2XL U81 ( .A(n85), .B(n100), .Y(n404) );
  NAND2XL U82 ( .A(n25), .B(n15), .Y(n339) );
  NAND2XL U83 ( .A(n97), .B(n20), .Y(n394) );
  NAND2XL U84 ( .A(n15), .B(n95), .Y(n458) );
  NAND2XL U85 ( .A(n81), .B(n247), .Y(n250) );
  NAND2XL U86 ( .A(n99), .B(n15), .Y(n362) );
  NAND2XL U87 ( .A(n85), .B(a[7]), .Y(n385) );
  NAND2XL U88 ( .A(n97), .B(n83), .Y(n466) );
  AOI22XL U89 ( .A0(n96), .A1(n431), .B0(n22), .B1(n430), .Y(n433) );
  INVXL U90 ( .A(n85), .Y(n224) );
  NAND2XL U91 ( .A(n7), .B(n22), .Y(n299) );
  NAND2XL U92 ( .A(n15), .B(a[1]), .Y(n296) );
  INVXL U93 ( .A(n97), .Y(n483) );
  XOR2XL U94 ( .A(n191), .B(n216), .Y(n203) );
  XOR3X2 U95 ( .A(n301), .B(n39), .C(n300), .Y(c[7]) );
  XNOR2X1 U96 ( .A(n296), .B(n473), .Y(n39) );
  OAI2BB1X1 U97 ( .A0N(n84), .A1N(n181), .B0(n180), .Y(n182) );
  AOI22XL U98 ( .A0(n28), .A1(n478), .B0(n30), .B1(n477), .Y(n481) );
  AOI22XL U99 ( .A0(n34), .A1(n397), .B0(n37), .B1(n396), .Y(n400) );
  AOI22XL U100 ( .A0(n24), .A1(n447), .B0(n98), .B1(n446), .Y(n449) );
  AOI22XL U101 ( .A0(n30), .A1(n487), .B0(n31), .B1(n486), .Y(n488) );
  NAND2XL U102 ( .A(n17), .B(n33), .Y(n233) );
  NAND2XL U103 ( .A(n99), .B(n87), .Y(n436) );
  NAND2BXL U104 ( .AN(b[2]), .B(n102), .Y(n141) );
  NAND2XL U105 ( .A(n86), .B(n100), .Y(n384) );
  NAND2XL U106 ( .A(n11), .B(n97), .Y(n149) );
  NAND2XL U107 ( .A(a[3]), .B(n92), .Y(n148) );
  NAND2BXL U108 ( .AN(n85), .B(n37), .Y(n226) );
  NOR2X1 U109 ( .A(n228), .B(n227), .Y(n236) );
  NAND2BXL U110 ( .AN(n85), .B(n36), .Y(n211) );
  NAND2XL U111 ( .A(n36), .B(n12), .Y(n359) );
  NAND2XL U112 ( .A(n34), .B(n87), .Y(n40) );
  XNOR2X1 U113 ( .A(n286), .B(n278), .Y(n43) );
  NAND2XL U114 ( .A(n28), .B(n92), .Y(n230) );
  NAND2XL U115 ( .A(n98), .B(n87), .Y(n427) );
  NAND2XL U116 ( .A(n84), .B(a[3]), .Y(n319) );
  NAND2XL U117 ( .A(n85), .B(a[8]), .Y(n69) );
  NAND2XL U118 ( .A(n101), .B(n84), .Y(n72) );
  NAND2XL U119 ( .A(b[9]), .B(n101), .Y(n234) );
  NAND2XL U120 ( .A(n100), .B(n87), .Y(n437) );
  NAND2XL U121 ( .A(n82), .B(n30), .Y(n402) );
  NAND2XL U122 ( .A(n99), .B(n12), .Y(n204) );
  INVXL U123 ( .A(n86), .Y(n382) );
  NAND2XL U124 ( .A(n101), .B(n92), .Y(n278) );
  NAND2XL U125 ( .A(n30), .B(n21), .Y(n254) );
  NAND2XL U126 ( .A(n100), .B(n11), .Y(n222) );
  NAND2XL U127 ( .A(a[7]), .B(n18), .Y(n435) );
  NAND2XL U128 ( .A(a[7]), .B(n87), .Y(n451) );
  NAND2X1 U129 ( .A(a[7]), .B(b[9]), .Y(n438) );
  XOR3X2 U130 ( .A(n47), .B(n316), .C(n315), .Y(n378) );
  NAND2XL U131 ( .A(n34), .B(n21), .Y(n47) );
  NAND2XL U132 ( .A(n18), .B(n22), .Y(n343) );
  NAND2XL U133 ( .A(n86), .B(n33), .Y(n205) );
  NAND2XL U134 ( .A(n100), .B(n92), .Y(n450) );
  NAND2XL U135 ( .A(n98), .B(n86), .Y(n358) );
  NAND2XL U136 ( .A(n30), .B(n11), .Y(n286) );
  AND2X1 U137 ( .A(n8), .B(n96), .Y(n79) );
  NAND2XL U138 ( .A(a[8]), .B(n87), .Y(n223) );
  NAND2XL U139 ( .A(n96), .B(n9), .Y(n363) );
  NAND2BXL U140 ( .AN(n86), .B(n37), .Y(n247) );
  NAND2XL U141 ( .A(n95), .B(n21), .Y(n365) );
  NAND2XL U142 ( .A(n24), .B(n18), .Y(n395) );
  NAND2XL U143 ( .A(n86), .B(a[7]), .Y(n426) );
  XNOR3X2 U144 ( .A(n49), .B(n50), .C(n214), .Y(n215) );
  NAND2XL U145 ( .A(b[9]), .B(n30), .Y(n49) );
  NAND2XL U146 ( .A(n17), .B(n101), .Y(n50) );
  AOI22XL U147 ( .A0(n34), .A1(n390), .B0(n31), .B1(n389), .Y(n391) );
  NAND2XL U148 ( .A(n82), .B(n31), .Y(n408) );
  NAND2XL U149 ( .A(n83), .B(n30), .Y(n407) );
  NAND2XL U150 ( .A(n8), .B(n24), .Y(n349) );
  NAND2XL U151 ( .A(a[3]), .B(n82), .Y(n467) );
  NAND2XL U152 ( .A(n95), .B(n12), .Y(n413) );
  INVXL U153 ( .A(n292), .Y(n221) );
  XOR3X2 U154 ( .A(n51), .B(n347), .C(n346), .Y(n351) );
  NAND2XL U155 ( .A(n30), .B(b[2]), .Y(n51) );
  NAND2XL U156 ( .A(n12), .B(n96), .Y(n133) );
  NAND2XL U157 ( .A(n92), .B(n97), .Y(n134) );
  NAND2XL U158 ( .A(n15), .B(n24), .Y(n331) );
  NAND2XL U159 ( .A(n8), .B(n97), .Y(n332) );
  NAND2XL U160 ( .A(n101), .B(n83), .Y(n68) );
  XOR2X1 U161 ( .A(n52), .B(n53), .Y(n412) );
  XNOR3X2 U162 ( .A(n403), .B(n372), .C(n371), .Y(n52) );
  XNOR2X1 U163 ( .A(n405), .B(n404), .Y(n53) );
  XOR2X1 U164 ( .A(n261), .B(n260), .Y(n266) );
  NAND2XL U165 ( .A(n28), .B(n12), .Y(n259) );
  AOI22XL U166 ( .A0(n97), .A1(n443), .B0(n24), .B1(n442), .Y(n445) );
  NAND2XL U167 ( .A(n100), .B(n18), .Y(n425) );
  NAND2XL U168 ( .A(n98), .B(n11), .Y(n439) );
  NAND2XL U169 ( .A(n99), .B(n92), .Y(n440) );
  INVXL U170 ( .A(n101), .Y(n398) );
  AND2X1 U171 ( .A(n98), .B(n92), .Y(n66) );
  OAI2BB1X1 U172 ( .A0N(n102), .A1N(n303), .B0(n374), .Y(n106) );
  AND2X1 U173 ( .A(n101), .B(n87), .Y(n253) );
  INVXL U174 ( .A(n37), .Y(n373) );
  INVXL U175 ( .A(n92), .Y(n109) );
  NAND2XL U176 ( .A(n18), .B(a[1]), .Y(n335) );
  NAND2XL U177 ( .A(n24), .B(n20), .Y(n415) );
  NAND2XL U178 ( .A(n96), .B(n21), .Y(n417) );
  NAND2XL U179 ( .A(n24), .B(b[2]), .Y(n455) );
  NAND2XL U180 ( .A(n22), .B(n9), .Y(n418) );
  NAND2XL U181 ( .A(n95), .B(n18), .Y(n317) );
  NAND2XL U182 ( .A(n25), .B(n18), .Y(n416) );
  NAND2XL U183 ( .A(n95), .B(n8), .Y(n297) );
  NAND2XL U184 ( .A(n24), .B(n6), .Y(n475) );
  NAND2BXL U185 ( .AN(b[1]), .B(n102), .Y(n126) );
  NAND2XL U186 ( .A(n81), .B(n126), .Y(n129) );
  NAND2XL U187 ( .A(b[0]), .B(n484), .Y(n55) );
  XNOR2X1 U188 ( .A(n140), .B(n361), .Y(n356) );
  XNOR2X1 U189 ( .A(n140), .B(n372), .Y(n195) );
  XNOR2X1 U190 ( .A(n216), .B(n58), .Y(n292) );
  XNOR2X1 U191 ( .A(n58), .B(n2), .Y(n324) );
  XNOR3X2 U192 ( .A(n173), .B(n170), .C(n169), .Y(n263) );
  XOR2X1 U193 ( .A(n434), .B(n435), .Y(n173) );
  XOR3X2 U194 ( .A(n154), .B(n436), .C(n66), .Y(n170) );
  XOR3X2 U195 ( .A(n168), .B(n167), .C(n166), .Y(n169) );
  INVX1 U196 ( .A(n192), .Y(n361) );
  XOR2X1 U197 ( .A(n266), .B(n3), .Y(n357) );
  INVX1 U198 ( .A(n359), .Y(n372) );
  NOR2X1 U199 ( .A(n380), .B(n382), .Y(n403) );
  XOR3X2 U200 ( .A(n63), .B(n338), .C(n337), .Y(c[9]) );
  XNOR3X2 U201 ( .A(n371), .B(n327), .C(n326), .Y(n338) );
  XNOR3X2 U202 ( .A(n336), .B(n335), .C(n334), .Y(n337) );
  XOR2X1 U203 ( .A(n325), .B(n489), .Y(n326) );
  XOR3X2 U204 ( .A(n357), .B(n356), .C(n355), .Y(c[10]) );
  XNOR3X2 U205 ( .A(n354), .B(n353), .C(n352), .Y(n355) );
  XNOR2X1 U206 ( .A(n343), .B(n339), .Y(n353) );
  XOR2X1 U207 ( .A(n351), .B(n350), .Y(n352) );
  XNOR3X2 U208 ( .A(n61), .B(n370), .C(n369), .Y(c[11]) );
  XOR3X2 U209 ( .A(n368), .B(n367), .C(n366), .Y(n369) );
  XNOR3X2 U210 ( .A(n400), .B(n361), .C(n360), .Y(n370) );
  XOR2X1 U211 ( .A(n364), .B(n394), .Y(n367) );
  XNOR3X2 U212 ( .A(n474), .B(n299), .C(n298), .Y(n300) );
  XOR2X1 U213 ( .A(n357), .B(n292), .Y(n301) );
  XOR2X1 U214 ( .A(n223), .B(n222), .Y(n237) );
  XOR3X2 U215 ( .A(n234), .B(n233), .C(n230), .Y(n235) );
  INVX1 U216 ( .A(n378), .Y(n330) );
  XNOR3X2 U217 ( .A(n361), .B(n193), .C(n174), .Y(n57) );
  XOR3X2 U218 ( .A(n59), .B(n60), .C(n215), .Y(n58) );
  XNOR2X1 U219 ( .A(n205), .B(n204), .Y(n59) );
  XOR2X1 U220 ( .A(n450), .B(n451), .Y(n60) );
  XOR2X1 U221 ( .A(n3), .B(n330), .Y(n61) );
  INVX1 U222 ( .A(n81), .Y(n304) );
  XNOR3X2 U223 ( .A(n195), .B(n174), .C(n191), .Y(n62) );
  XNOR3X2 U224 ( .A(n324), .B(n57), .C(n246), .Y(c[5]) );
  XNOR3X2 U225 ( .A(n454), .B(n240), .C(n239), .Y(n246) );
  XOR2X1 U226 ( .A(n238), .B(n455), .Y(n239) );
  XNOR3X2 U227 ( .A(n324), .B(n61), .C(n323), .Y(c[8]) );
  XOR3X2 U228 ( .A(n481), .B(n322), .C(n321), .Y(n323) );
  XOR3X2 U229 ( .A(n482), .B(n79), .C(n320), .Y(n321) );
  XNOR3X2 U230 ( .A(n203), .B(n202), .C(n196), .Y(c[3]) );
  XNOR3X2 U231 ( .A(n441), .B(n195), .C(n194), .Y(n196) );
  XOR2X1 U232 ( .A(n193), .B(n192), .Y(n202) );
  XNOR2X1 U233 ( .A(n266), .B(n2), .Y(n63) );
  NOR2XL U234 ( .A(n480), .B(n380), .Y(n473) );
  NOR2BX1 U235 ( .AN(n103), .B(n92), .Y(n104) );
  XNOR2X1 U236 ( .A(n445), .B(n444), .Y(n194) );
  OAI2BB1X1 U237 ( .A0N(n12), .A1N(n122), .B0(n111), .Y(n192) );
  OAI21XL U238 ( .A0(n30), .A1(n35), .B0(n38), .Y(n478) );
  OAI21XL U239 ( .A0(n28), .A1(n485), .B0(n5), .Y(n477) );
  OAI21XL U240 ( .A0(n13), .A1(n35), .B0(n38), .Y(n453) );
  OAI21XL U241 ( .A0(n98), .A1(n485), .B0(n55), .Y(n452) );
  OAI21XL U242 ( .A0(n37), .A1(n35), .B0(n38), .Y(n397) );
  OAI21XL U243 ( .A0(n34), .A1(n485), .B0(n55), .Y(n396) );
  AOI22X1 U244 ( .A0(n26), .A1(n472), .B0(n28), .B1(n471), .Y(n474) );
  OAI21XL U245 ( .A0(n28), .A1(n35), .B0(n38), .Y(n472) );
  OAI21XL U246 ( .A0(n26), .A1(n14), .B0(n55), .Y(n471) );
  OAI21XL U247 ( .A0(n98), .A1(n35), .B0(n38), .Y(n447) );
  OAI21XL U248 ( .A0(n24), .A1(n485), .B0(n5), .Y(n446) );
  AOI21X1 U249 ( .A0(n81), .A1(n226), .B0(n382), .Y(n227) );
  OAI21XL U250 ( .A0(n100), .A1(n484), .B0(n54), .Y(n462) );
  OAI21XL U251 ( .A0(n24), .A1(n35), .B0(n38), .Y(n443) );
  OAI21XL U252 ( .A0(n22), .A1(n35), .B0(n38), .Y(n431) );
  OAI21XL U253 ( .A0(n31), .A1(n485), .B0(n5), .Y(n390) );
  OAI21XL U254 ( .A0(n34), .A1(n35), .B0(n38), .Y(n389) );
  OAI21XL U255 ( .A0(n99), .A1(n485), .B0(n5), .Y(n461) );
  OAI21XL U256 ( .A0(n97), .A1(n485), .B0(n55), .Y(n442) );
  OAI21XL U257 ( .A0(n96), .A1(n14), .B0(n5), .Y(n430) );
  OAI2BB1X2 U258 ( .A0N(n92), .A1N(n106), .B0(n105), .Y(n108) );
  XNOR3X2 U259 ( .A(n427), .B(n151), .C(n150), .Y(n152) );
  XNOR3X2 U260 ( .A(n147), .B(n146), .C(n145), .Y(n153) );
  INVX1 U261 ( .A(b[2]), .Y(n480) );
  OAI21XL U262 ( .A0(n305), .A1(n304), .B0(n9), .Y(n306) );
  NOR2BX1 U263 ( .AN(n37), .B(n20), .Y(n305) );
  OAI2BB1X1 U264 ( .A0N(n82), .A1N(n144), .B0(n143), .Y(n146) );
  NAND2X1 U265 ( .A(n101), .B(n12), .Y(n316) );
  OAI2BB1X1 U266 ( .A0N(n20), .A1N(n314), .B0(n306), .Y(n315) );
  XOR2X1 U267 ( .A(n259), .B(n254), .Y(n260) );
  XNOR3X2 U268 ( .A(n253), .B(n252), .C(n251), .Y(n261) );
  XNOR3X2 U269 ( .A(n437), .B(n438), .C(n175), .Y(n190) );
  XNOR3X2 U270 ( .A(n188), .B(n187), .C(n182), .Y(n189) );
  NAND2X1 U271 ( .A(n20), .B(n34), .Y(n252) );
  XOR2X1 U272 ( .A(n139), .B(n138), .Y(n191) );
  XNOR3X2 U273 ( .A(n384), .B(n137), .C(n136), .Y(n138) );
  XNOR3X2 U274 ( .A(n132), .B(n131), .C(n130), .Y(n139) );
  XNOR3X2 U275 ( .A(n64), .B(n65), .C(n317), .Y(n322) );
  OR2X2 U276 ( .A(n480), .B(n479), .Y(n64) );
  OAI2BB1X1 U277 ( .A0N(n20), .A1N(n290), .B0(n289), .Y(n291) );
  XOR2X1 U278 ( .A(n162), .B(n155), .Y(n167) );
  XOR2X1 U279 ( .A(n149), .B(n148), .Y(n151) );
  NAND2X1 U280 ( .A(n17), .B(a[8]), .Y(n177) );
  XOR2X1 U281 ( .A(n386), .B(n387), .Y(n137) );
  NAND2X1 U282 ( .A(n98), .B(b[9]), .Y(n386) );
  XOR3X2 U283 ( .A(n413), .B(n414), .C(n378), .Y(n422) );
  XOR2X1 U284 ( .A(n412), .B(n411), .Y(n414) );
  XOR2X1 U285 ( .A(n410), .B(n409), .Y(n411) );
  XNOR3X2 U286 ( .A(n62), .B(n221), .C(n220), .Y(c[4]) );
  XNOR3X2 U287 ( .A(n449), .B(n219), .C(n218), .Y(n220) );
  NAND2X1 U288 ( .A(a[0]), .B(n6), .Y(n219) );
  NAND2X1 U289 ( .A(n95), .B(n9), .Y(n346) );
  NAND2X1 U290 ( .A(n20), .B(n96), .Y(n347) );
  XOR2X1 U291 ( .A(n408), .B(n407), .Y(n409) );
  XOR2X1 U292 ( .A(n467), .B(n466), .Y(n468) );
  XOR3X2 U293 ( .A(n393), .B(n392), .C(n391), .Y(n354) );
  NAND2X1 U294 ( .A(n83), .B(n26), .Y(n392) );
  NAND2X1 U295 ( .A(b[3]), .B(n28), .Y(n393) );
  OAI2BB1X1 U296 ( .A0N(n37), .A1N(n210), .B0(n81), .Y(n213) );
  NAND2X1 U297 ( .A(n100), .B(n20), .Y(n434) );
  OAI2BB1X1 U298 ( .A0N(n82), .A1N(n165), .B0(n164), .Y(n166) );
  OAI21XL U299 ( .A0(n163), .A1(n304), .B0(n83), .Y(n164) );
  NOR2BX1 U300 ( .AN(n102), .B(n82), .Y(n163) );
  XNOR3X2 U301 ( .A(n67), .B(n68), .C(n385), .Y(n130) );
  XOR3X2 U302 ( .A(n135), .B(n134), .C(n133), .Y(n136) );
  NOR2BX1 U303 ( .AN(n103), .B(n84), .Y(n179) );
  OAI2BB1X1 U304 ( .A0N(n18), .A1N(n250), .B0(n249), .Y(n251) );
  AOI21X1 U305 ( .A0(n85), .A1(n213), .B0(n212), .Y(n214) );
  XOR2X1 U306 ( .A(n465), .B(n464), .Y(n469) );
  NOR2X1 U307 ( .A(n480), .B(n463), .Y(n464) );
  INVX1 U308 ( .A(n98), .Y(n463) );
  XOR2X1 U309 ( .A(n377), .B(n406), .Y(n410) );
  NAND2X1 U310 ( .A(b[2]), .B(n34), .Y(n406) );
  NAND2X1 U311 ( .A(n84), .B(n28), .Y(n405) );
  XOR2X1 U312 ( .A(n470), .B(n460), .Y(n265) );
  XOR2X1 U313 ( .A(n459), .B(n458), .Y(n460) );
  XOR2X1 U314 ( .A(n469), .B(n468), .Y(n470) );
  NAND2X1 U315 ( .A(n84), .B(n96), .Y(n459) );
  NOR2BX1 U316 ( .AN(n103), .B(n82), .Y(n142) );
  NOR2BX1 U317 ( .AN(n36), .B(n20), .Y(n288) );
  NOR2BX1 U318 ( .AN(n103), .B(n17), .Y(n248) );
  NOR2BX1 U319 ( .AN(n36), .B(n12), .Y(n110) );
  NOR2BX1 U320 ( .AN(n103), .B(b[2]), .Y(n127) );
  XOR2X1 U321 ( .A(n330), .B(n488), .Y(n336) );
  OAI21XL U322 ( .A0(n31), .A1(n35), .B0(n38), .Y(n487) );
  OAI21XL U323 ( .A0(n30), .A1(n485), .B0(n55), .Y(n486) );
  NAND2BXL U324 ( .AN(n86), .B(n103), .Y(n225) );
  AND2X2 U325 ( .A(n12), .B(a[3]), .Y(n154) );
  XNOR3X2 U326 ( .A(n69), .B(n72), .C(n426), .Y(n145) );
  AND2X2 U327 ( .A(n33), .B(n82), .Y(n132) );
  AND2X2 U328 ( .A(n34), .B(n83), .Y(n147) );
  AND2X2 U329 ( .A(n34), .B(n84), .Y(n168) );
  XNOR2X1 U330 ( .A(n428), .B(n425), .Y(n150) );
  NOR2X1 U331 ( .A(n381), .B(n480), .Y(n432) );
  XOR2X1 U332 ( .A(n439), .B(n440), .Y(n175) );
  INVX1 U333 ( .A(n100), .Y(n479) );
  INVX1 U334 ( .A(n84), .Y(n210) );
  INVX1 U335 ( .A(n87), .Y(n303) );
  INVX1 U336 ( .A(n83), .Y(n178) );
  AOI22X1 U337 ( .A0(a[0]), .A1(n424), .B0(a[1]), .B1(n423), .Y(n429) );
  OAI21XL U338 ( .A0(a[1]), .A1(n35), .B0(n38), .Y(n424) );
  OAI21XL U339 ( .A0(n95), .A1(n14), .B0(n5), .Y(n423) );
  XNOR2X1 U340 ( .A(n457), .B(n456), .Y(n240) );
  NAND2X1 U341 ( .A(n6), .B(n96), .Y(n456) );
  NOR2X1 U342 ( .A(n381), .B(n14), .Y(n388) );
  XOR3X2 U343 ( .A(n399), .B(n395), .C(n365), .Y(n366) );
  NOR2X1 U344 ( .A(n398), .B(n480), .Y(n399) );
  NOR2X1 U345 ( .A(n381), .B(n383), .Y(n441) );
  INVX1 U346 ( .A(n82), .Y(n383) );
  XNOR2X1 U347 ( .A(n77), .B(n78), .Y(n327) );
  AND2X2 U348 ( .A(b[3]), .B(n26), .Y(n77) );
  NAND2X1 U349 ( .A(n28), .B(b[2]), .Y(n78) );
  XOR2X1 U350 ( .A(n349), .B(n348), .Y(n350) );
  XOR2X1 U351 ( .A(n420), .B(n419), .Y(n421) );
  XOR2X1 U352 ( .A(n416), .B(n415), .Y(n420) );
  XOR2X1 U353 ( .A(n418), .B(n417), .Y(n419) );
  NAND2X1 U354 ( .A(n95), .B(n7), .Y(n238) );
  NAND2X1 U355 ( .A(n26), .B(n7), .Y(n364) );
  NAND2X1 U356 ( .A(n25), .B(n7), .Y(n325) );
  XNOR2X1 U357 ( .A(n319), .B(n318), .Y(n320) );
  XOR3X2 U358 ( .A(n333), .B(n332), .C(n331), .Y(n334) );
  NAND2X1 U359 ( .A(n95), .B(n20), .Y(n333) );
  XOR3X2 U360 ( .A(n476), .B(n475), .C(n297), .Y(n298) );
  NAND2X1 U361 ( .A(n25), .B(b[3]), .Y(n476) );
  NAND2X1 U362 ( .A(n98), .B(n83), .Y(n482) );
  INVX1 U363 ( .A(n95), .Y(n381) );
  XOR2X1 U364 ( .A(n363), .B(n362), .Y(n368) );
  XNOR3X2 U365 ( .A(n359), .B(n401), .C(n80), .Y(n360) );
  XNOR2X1 U366 ( .A(n358), .B(n402), .Y(n80) );
  NAND2X1 U367 ( .A(n83), .B(n28), .Y(n401) );
  XOR2X1 U368 ( .A(n217), .B(n448), .Y(n218) );
  NAND2X1 U369 ( .A(b[3]), .B(a[1]), .Y(n217) );
  NOR2X1 U370 ( .A(n480), .B(n483), .Y(n448) );
  INVX1 U371 ( .A(b[0]), .Y(n485) );
  INVX1 U372 ( .A(b[1]), .Y(n484) );
  OAI2BB1X1 U373 ( .A0N(b[2]), .A1N(n129), .B0(n128), .Y(n131) );
  BUFX3 U374 ( .A(a[4]), .Y(n98) );
  BUFX3 U375 ( .A(a[6]), .Y(n100) );
  BUFX3 U376 ( .A(a[1]), .Y(n96) );
  XOR2X1 U377 ( .A(n422), .B(n421), .Y(c[12]) );
  BUFX3 U378 ( .A(a[9]), .Y(n101) );
  BUFX3 U379 ( .A(b[3]), .Y(n82) );
  BUFX3 U380 ( .A(b[11]), .Y(n92) );
  BUFX3 U381 ( .A(b[6]), .Y(n85) );
  BUFX3 U382 ( .A(b[10]), .Y(n87) );
  BUFX3 U383 ( .A(b[7]), .Y(n86) );
  BUFX3 U384 ( .A(b[4]), .Y(n83) );
  BUFX3 U385 ( .A(b[5]), .Y(n84) );
  XNOR3X2 U386 ( .A(n63), .B(n265), .C(n264), .Y(c[6]) );
  XNOR2X1 U387 ( .A(n57), .B(n4), .Y(c[2]) );
  XNOR3X2 U388 ( .A(n388), .B(n356), .C(n191), .Y(c[0]) );
  BUFX3 U389 ( .A(a[0]), .Y(n95) );
  OAI21XL U390 ( .A0(n110), .A1(n375), .B0(n21), .Y(n111) );
  OAI21XL U391 ( .A0(n288), .A1(n375), .B0(n18), .Y(n289) );
  OAI21XL U392 ( .A0(n127), .A1(n375), .B0(b[1]), .Y(n128) );
  AOI21XL U393 ( .A0(n302), .A1(n225), .B0(n224), .Y(n228) );
  AOI2BB2X1 U394 ( .B0(b[0]), .B1(n375), .A0N(n81), .A1N(n484), .Y(n376) );
  OAI21XL U395 ( .A0(n248), .A1(n375), .B0(n86), .Y(n249) );
  OAI21XL U396 ( .A0(n142), .A1(n375), .B0(b[2]), .Y(n143) );
  OAI2BB1X1 U397 ( .A0N(n103), .A1N(n178), .B0(n302), .Y(n165) );
  AOI21X1 U398 ( .A0(n302), .A1(n211), .B0(n210), .Y(n212) );
  OAI21XL U399 ( .A0(n179), .A1(n375), .B0(n83), .Y(n180) );
  XOR2X4 U400 ( .A(n108), .B(n107), .Y(n371) );
endmodule


module multiplier_0 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n36, n37, n38, n39, n43, n47, n50, n51, n52, n53,
         n54, n55, n57, n58, n59, n61, n62, n63, n64, n77, n81, n83, n84, n85,
         n86, n87, n92, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n122, n126, n127, n128,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n162, n163, n164, n165, n166, n167, n168, n169, n170, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n187, n189,
         n192, n193, n194, n195, n202, n203, n204, n205, n210, n211, n212,
         n213, n214, n215, n216, n217, n219, n220, n221, n225, n239, n240,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n259, n260,
         n261, n262, n263, n264, n265, n266, n286, n288, n289, n290, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n311, n314, n315, n316, n317, n318, n319, n320, n321, n323, n324,
         n325, n326, n327, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n380, n381, n385, n386, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559;

  AOI21X2 U1 ( .A0(n98), .A1(n127), .B0(n126), .Y(n128) );
  INVX1 U2 ( .A(n357), .Y(n367) );
  BUFX4 U3 ( .A(a[12]), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n13), .A1N(n38), .B0(n368), .Y(n212) );
  OAI211X1 U5 ( .A0(n400), .A1(n357), .B0(n369), .C0(n368), .Y(n370) );
  NOR2X1 U6 ( .A(n23), .B(n39), .Y(n264) );
  NAND2BX2 U7 ( .AN(n109), .B(n110), .Y(n357) );
  NAND2BX1 U8 ( .AN(n483), .B(n482), .Y(n52) );
  NOR2XL U9 ( .A(n34), .B(n47), .Y(n289) );
  NOR2X1 U10 ( .A(n367), .B(n540), .Y(n358) );
  NOR2X1 U11 ( .A(n50), .B(n39), .Y(n303) );
  NAND2BX1 U12 ( .AN(n482), .B(n483), .Y(n51) );
  XOR3X2 U13 ( .A(n321), .B(n320), .C(n556), .Y(n323) );
  NAND2X1 U14 ( .A(n51), .B(n52), .Y(n2) );
  XNOR3X2 U15 ( .A(n151), .B(n356), .C(n432), .Y(n86) );
  OAI221XL U16 ( .A0(n361), .A1(n111), .B0(n64), .B1(n39), .C0(n365), .Y(n366)
         );
  XOR3X2 U17 ( .A(n408), .B(n407), .C(n415), .Y(n416) );
  XOR3X2 U18 ( .A(n2), .B(n151), .C(n402), .Y(n496) );
  XOR3X2 U19 ( .A(n473), .B(n472), .C(n480), .Y(n483) );
  OAI2BB1X1 U20 ( .A0N(n17), .A1N(n109), .B0(n368), .Y(n182) );
  NOR2X1 U21 ( .A(n7), .B(n540), .Y(n431) );
  XNOR3X2 U22 ( .A(n497), .B(n496), .C(n495), .Y(c[3]) );
  XOR2X1 U23 ( .A(n468), .B(n469), .Y(n473) );
  OAI2BB1X1 U24 ( .A0N(n4), .A1N(n371), .B0(n370), .Y(n468) );
  AND2X2 U25 ( .A(n51), .B(n52), .Y(n1) );
  AOI21X1 U26 ( .A0(n363), .A1(n122), .B0(n47), .Y(n131) );
  XOR2X1 U27 ( .A(n143), .B(n142), .Y(n145) );
  XOR2X1 U28 ( .A(n402), .B(n57), .Y(n438) );
  INVX1 U29 ( .A(n320), .Y(n325) );
  XOR2X1 U30 ( .A(n503), .B(n176), .Y(n193) );
  INVX1 U31 ( .A(n151), .Y(n373) );
  XNOR3X2 U32 ( .A(n61), .B(n77), .C(n402), .Y(n81) );
  XNOR3X2 U33 ( .A(n289), .B(n288), .C(n286), .Y(n3) );
  INVX1 U34 ( .A(n377), .Y(n495) );
  INVX1 U35 ( .A(b[10]), .Y(n47) );
  INVX1 U36 ( .A(b[4]), .Y(n4) );
  INVX1 U37 ( .A(n4), .Y(n5) );
  BUFX3 U38 ( .A(b[3]), .Y(n6) );
  BUFX3 U39 ( .A(b[3]), .Y(n99) );
  INVX1 U40 ( .A(a[9]), .Y(n7) );
  INVX1 U41 ( .A(n7), .Y(n8) );
  INVX1 U42 ( .A(n7), .Y(n9) );
  BUFX3 U43 ( .A(n64), .Y(n10) );
  INVX1 U44 ( .A(n385), .Y(n11) );
  INVX1 U45 ( .A(n101), .Y(n385) );
  INVX1 U46 ( .A(b[1]), .Y(n12) );
  INVX1 U47 ( .A(b[7]), .Y(n13) );
  INVX1 U48 ( .A(n13), .Y(n14) );
  CLKINVX2 U49 ( .A(n13), .Y(n15) );
  NAND2X1 U50 ( .A(n14), .B(n8), .Y(n163) );
  INVX1 U51 ( .A(n378), .Y(n16) );
  INVX1 U52 ( .A(b[5]), .Y(n17) );
  INVX1 U53 ( .A(n17), .Y(n18) );
  INVX1 U54 ( .A(n17), .Y(n19) );
  INVX1 U55 ( .A(b[8]), .Y(n20) );
  INVXL U56 ( .A(n20), .Y(n21) );
  INVX1 U57 ( .A(b[9]), .Y(n22) );
  INVXL U58 ( .A(n22), .Y(n23) );
  BUFX3 U59 ( .A(b[11]), .Y(n24) );
  INVX1 U60 ( .A(n550), .Y(n25) );
  INVX1 U61 ( .A(n481), .Y(n26) );
  INVX1 U62 ( .A(n519), .Y(n27) );
  INVX1 U63 ( .A(n539), .Y(n28) );
  INVX1 U64 ( .A(a[7]), .Y(n29) );
  INVX1 U65 ( .A(n29), .Y(n30) );
  INVX1 U66 ( .A(a[8]), .Y(n31) );
  INVX1 U67 ( .A(n31), .Y(n32) );
  INVX1 U68 ( .A(n31), .Y(n33) );
  INVX1 U69 ( .A(a[10]), .Y(n34) );
  INVX1 U70 ( .A(n34), .Y(n36) );
  INVX1 U71 ( .A(n34), .Y(n37) );
  AND2X2 U72 ( .A(n37), .B(n101), .Y(n132) );
  BUFX3 U73 ( .A(n109), .Y(n38) );
  CLKBUFX8 U74 ( .A(a[11]), .Y(n109) );
  INVX1 U75 ( .A(n110), .Y(n39) );
  INVX1 U76 ( .A(n39), .Y(n43) );
  NAND2X1 U77 ( .A(b[0]), .B(n552), .Y(n64) );
  XNOR3X4 U78 ( .A(n53), .B(n376), .C(n375), .Y(n512) );
  XNOR3X4 U79 ( .A(n533), .B(n53), .C(n58), .Y(n401) );
  XOR3X4 U80 ( .A(n54), .B(n253), .C(n252), .Y(n53) );
  AND2X2 U81 ( .A(n15), .B(n36), .Y(n176) );
  NOR2X2 U82 ( .A(n248), .B(n247), .Y(n253) );
  AOI21XL U83 ( .A0(n363), .A1(n240), .B0(n239), .Y(n248) );
  AOI21XL U84 ( .A0(n98), .A1(n246), .B0(n386), .Y(n247) );
  XOR2X2 U85 ( .A(n372), .B(n58), .Y(n290) );
  XNOR3X4 U86 ( .A(n193), .B(n192), .C(n189), .Y(n58) );
  OAI2BB1XL U87 ( .A0N(n43), .A1N(n385), .B0(n363), .Y(n150) );
  XNOR2X4 U88 ( .A(n133), .B(n132), .Y(n320) );
  XNOR2X1 U89 ( .A(n260), .B(n53), .Y(n84) );
  XNOR2X4 U90 ( .A(n320), .B(n355), .Y(n402) );
  XOR2X2 U91 ( .A(n164), .B(n163), .Y(n170) );
  AOI21X1 U92 ( .A0(n400), .A1(n109), .B0(n4), .Y(n369) );
  XOR2X4 U93 ( .A(n548), .B(n547), .Y(n549) );
  XOR2X4 U94 ( .A(n401), .B(n536), .Y(n548) );
  NAND2XL U95 ( .A(b[1]), .B(n553), .Y(n551) );
  INVX1 U96 ( .A(n47), .Y(n50) );
  NAND2XL U97 ( .A(n105), .B(n50), .Y(n418) );
  NAND2XL U98 ( .A(n107), .B(b[10]), .Y(n477) );
  NAND2XL U99 ( .A(n32), .B(b[10]), .Y(n225) );
  NAND2BX1 U100 ( .AN(n109), .B(n110), .Y(n363) );
  NOR2X1 U101 ( .A(n385), .B(n481), .Y(n482) );
  BUFX3 U102 ( .A(b[6]), .Y(n100) );
  NAND2X1 U103 ( .A(b[9]), .B(n32), .Y(n179) );
  NOR2BX1 U104 ( .AN(n110), .B(b[8]), .Y(n210) );
  INVXL U105 ( .A(n98), .Y(n364) );
  NOR2X2 U106 ( .A(n131), .B(n128), .Y(n133) );
  XOR3X2 U107 ( .A(n337), .B(n422), .C(n336), .Y(n338) );
  XOR3X2 U108 ( .A(n290), .B(n203), .C(n204), .Y(c[4]) );
  NAND2X1 U109 ( .A(b[8]), .B(n32), .Y(n164) );
  NAND2X1 U110 ( .A(n108), .B(b[9]), .Y(n474) );
  NAND2XL U111 ( .A(n104), .B(n24), .Y(n417) );
  NAND2XL U112 ( .A(n103), .B(n6), .Y(n202) );
  XNOR2X1 U113 ( .A(n225), .B(n221), .Y(n54) );
  INVX2 U114 ( .A(n363), .Y(n302) );
  NOR2XL U115 ( .A(n380), .B(n386), .Y(n533) );
  XOR3X2 U116 ( .A(n300), .B(n55), .C(n299), .Y(c[7]) );
  XOR2X1 U117 ( .A(n531), .B(n529), .Y(n55) );
  NOR2XL U118 ( .A(n378), .B(n386), .Y(n57) );
  XOR2X1 U119 ( .A(n260), .B(n3), .Y(n339) );
  NAND2XL U120 ( .A(n43), .B(n101), .Y(n355) );
  AOI22XL U121 ( .A0(n28), .A1(n528), .B0(n30), .B1(n527), .Y(n530) );
  AOI22XL U122 ( .A0(n26), .A1(n499), .B0(n106), .B1(n498), .Y(n501) );
  NAND2XL U123 ( .A(n16), .B(n19), .Y(n326) );
  NAND2XL U124 ( .A(n15), .B(n105), .Y(n327) );
  AOI22XL U125 ( .A0(n37), .A1(n421), .B0(n9), .B1(n420), .Y(n423) );
  AOI22XL U126 ( .A0(n107), .A1(n518), .B0(n108), .B1(n517), .Y(n521) );
  NAND2BXL U127 ( .AN(b[10]), .B(n109), .Y(n127) );
  NAND2XL U128 ( .A(n6), .B(n28), .Y(n558) );
  NAND2XL U129 ( .A(n21), .B(n25), .Y(n334) );
  NAND2XL U130 ( .A(b[9]), .B(n37), .Y(n214) );
  NAND2XL U131 ( .A(n107), .B(n101), .Y(n178) );
  NAND2XL U132 ( .A(n99), .B(n110), .Y(n371) );
  NAND2XL U133 ( .A(n15), .B(n32), .Y(n470) );
  NAND2XL U134 ( .A(n19), .B(n102), .Y(n92) );
  NAND2XL U135 ( .A(n105), .B(n6), .Y(n523) );
  NAND2XL U136 ( .A(n104), .B(n101), .Y(n143) );
  NAND2XL U137 ( .A(n105), .B(b[11]), .Y(n142) );
  NAND2XL U138 ( .A(n6), .B(n33), .Y(n434) );
  NAND2XL U139 ( .A(n5), .B(n30), .Y(n433) );
  INVXL U140 ( .A(n106), .Y(n519) );
  INVXL U141 ( .A(n15), .Y(n386) );
  NAND2BXL U142 ( .AN(n100), .B(n109), .Y(n246) );
  NAND2XL U143 ( .A(n98), .B(n263), .Y(n266) );
  NAND2BXL U144 ( .AN(n21), .B(n38), .Y(n263) );
  NAND2XL U145 ( .A(n18), .B(n36), .Y(n469) );
  NAND2XL U146 ( .A(n15), .B(a[7]), .Y(n460) );
  NAND2XL U147 ( .A(a[7]), .B(n23), .Y(n486) );
  XNOR3X2 U148 ( .A(n59), .B(n428), .C(n306), .Y(n559) );
  NAND2XL U149 ( .A(n9), .B(n101), .Y(n59) );
  NAND2XL U150 ( .A(n104), .B(n23), .Y(n426) );
  NAND2XL U151 ( .A(n5), .B(n16), .Y(n557) );
  AOI22XL U152 ( .A0(n33), .A1(n555), .B0(n9), .B1(n554), .Y(n556) );
  NAND2XL U153 ( .A(n102), .B(n23), .Y(n318) );
  NAND2XL U154 ( .A(n15), .B(n104), .Y(n317) );
  NAND2XL U155 ( .A(n108), .B(n50), .Y(n485) );
  NAND2XL U156 ( .A(n15), .B(n108), .Y(n409) );
  NAND2XL U157 ( .A(n6), .B(n30), .Y(n425) );
  NAND2XL U158 ( .A(n5), .B(n28), .Y(n424) );
  NAND2XL U159 ( .A(n108), .B(n19), .Y(n346) );
  NAND2XL U160 ( .A(b[6]), .B(n104), .Y(n534) );
  NAND2XL U161 ( .A(n5), .B(n33), .Y(n440) );
  XOR2X1 U162 ( .A(n418), .B(n417), .Y(n61) );
  NAND2XL U163 ( .A(n33), .B(n24), .Y(n216) );
  NAND2XL U164 ( .A(n9), .B(b[11]), .Y(n261) );
  NAND2XL U165 ( .A(n100), .B(n30), .Y(n410) );
  NAND2XL U166 ( .A(n6), .B(n9), .Y(n441) );
  INVXL U167 ( .A(n109), .Y(n361) );
  NAND2XL U168 ( .A(n105), .B(n21), .Y(n427) );
  NAND2XL U169 ( .A(n19), .B(n103), .Y(n515) );
  NAND2XL U170 ( .A(b[6]), .B(n102), .Y(n514) );
  INVXL U171 ( .A(n107), .Y(n378) );
  NAND2XL U172 ( .A(n107), .B(n100), .Y(n347) );
  NAND2XL U173 ( .A(n33), .B(n101), .Y(n262) );
  NAND2XL U174 ( .A(a[7]), .B(b[10]), .Y(n503) );
  NAND2XL U175 ( .A(n98), .B(n165), .Y(n168) );
  OAI21XL U176 ( .A0(n166), .A1(n302), .B0(n5), .Y(n167) );
  NAND2BXL U177 ( .AN(b[4]), .B(n38), .Y(n165) );
  NAND2XL U178 ( .A(n21), .B(n9), .Y(n177) );
  XOR2X1 U179 ( .A(n220), .B(n219), .Y(n260) );
  NAND2XL U180 ( .A(n30), .B(n101), .Y(n217) );
  NAND2XL U181 ( .A(b[6]), .B(n105), .Y(n314) );
  NAND2XL U182 ( .A(n103), .B(n21), .Y(n311) );
  NAND2XL U183 ( .A(n102), .B(n11), .Y(n446) );
  XOR2X1 U184 ( .A(n147), .B(n146), .Y(n152) );
  NAND2XL U185 ( .A(n106), .B(n50), .Y(n461) );
  NAND2XL U186 ( .A(a[7]), .B(b[8]), .Y(n475) );
  NAND2XL U187 ( .A(n19), .B(n30), .Y(n436) );
  NAND2XL U188 ( .A(n100), .B(n28), .Y(n435) );
  NAND2XL U189 ( .A(n107), .B(n21), .Y(n412) );
  NAND2XL U190 ( .A(n106), .B(n23), .Y(n411) );
  NAND2XL U191 ( .A(b[4]), .B(n9), .Y(n406) );
  NAND2XL U192 ( .A(n18), .B(n33), .Y(n405) );
  NAND2XL U193 ( .A(n107), .B(n6), .Y(n544) );
  NAND2XL U194 ( .A(n106), .B(n5), .Y(n543) );
  NAND2BXL U195 ( .AN(b[11]), .B(n110), .Y(n122) );
  XNOR3X2 U196 ( .A(n62), .B(n549), .C(n353), .Y(c[8]) );
  NAND2XL U197 ( .A(n21), .B(a[0]), .Y(n62) );
  NAND2XL U198 ( .A(n27), .B(b[6]), .Y(n330) );
  NAND2XL U199 ( .A(n102), .B(n50), .Y(n331) );
  NAND2XL U200 ( .A(n103), .B(n23), .Y(n332) );
  NAND2XL U201 ( .A(n103), .B(n50), .Y(n349) );
  NAND2XL U202 ( .A(n102), .B(n24), .Y(n350) );
  AOI22XL U203 ( .A0(n30), .A1(n538), .B0(n33), .B1(n537), .Y(n542) );
  INVXL U204 ( .A(n108), .Y(n539) );
  XNOR2X1 U205 ( .A(n63), .B(n83), .Y(c[0]) );
  XOR2X1 U206 ( .A(n377), .B(n419), .Y(n63) );
  NAND2XL U207 ( .A(n105), .B(n19), .Y(n535) );
  BUFX8 U208 ( .A(n368), .Y(n98) );
  NAND2XL U209 ( .A(n24), .B(n37), .Y(n428) );
  NAND2XL U210 ( .A(n107), .B(b[9]), .Y(n462) );
  NAND2XL U211 ( .A(n108), .B(b[8]), .Y(n459) );
  AOI22XL U212 ( .A0(n37), .A1(n430), .B0(n38), .B1(n429), .Y(n432) );
  NAND2XL U213 ( .A(n106), .B(n101), .Y(n487) );
  NAND2XL U214 ( .A(n107), .B(n24), .Y(n488) );
  OAI2BB1X1 U215 ( .A0N(n21), .A1N(n212), .B0(n211), .Y(n213) );
  OAI21XL U216 ( .A0(n210), .A1(n302), .B0(n15), .Y(n211) );
  XOR2X1 U217 ( .A(n187), .B(n502), .Y(n189) );
  NAND2XL U218 ( .A(n108), .B(n24), .Y(n502) );
  AND2X1 U219 ( .A(n8), .B(n50), .Y(n215) );
  AND2X1 U220 ( .A(b[4]), .B(n36), .Y(n141) );
  AND2X1 U221 ( .A(n100), .B(n36), .Y(n173) );
  AND2X1 U222 ( .A(n106), .B(n15), .Y(n354) );
  NAND2XL U223 ( .A(n98), .B(n301), .Y(n305) );
  NAND2BXL U224 ( .AN(n23), .B(n38), .Y(n301) );
  NAND2XL U225 ( .A(n32), .B(n100), .Y(n95) );
  XOR2X1 U226 ( .A(n471), .B(n470), .Y(n472) );
  NAND2XL U227 ( .A(n100), .B(n8), .Y(n471) );
  INVX1 U228 ( .A(n99), .Y(n400) );
  NAND2XL U229 ( .A(a[1]), .B(b[6]), .Y(n298) );
  NAND2XL U230 ( .A(n26), .B(n23), .Y(n449) );
  NAND2XL U231 ( .A(n5), .B(n103), .Y(n508) );
  NAND2XL U232 ( .A(n27), .B(n21), .Y(n450) );
  NAND2XL U233 ( .A(n25), .B(n6), .Y(n509) );
  NAND2XL U234 ( .A(n26), .B(n5), .Y(n531) );
  NAND2XL U235 ( .A(n25), .B(n50), .Y(n452) );
  NAND2XL U236 ( .A(n103), .B(n24), .Y(n451) );
  NAND2XL U237 ( .A(n102), .B(n15), .Y(n295) );
  NAND2XL U238 ( .A(n19), .B(n25), .Y(n296) );
  NAND2XL U239 ( .A(n27), .B(n6), .Y(n532) );
  INVXL U240 ( .A(b[2]), .Y(n540) );
  NAND2XL U241 ( .A(n30), .B(b[2]), .Y(n96) );
  NAND2XL U242 ( .A(n106), .B(n19), .Y(n97) );
  OAI2BB1X1 U243 ( .A0N(n99), .A1N(n137), .B0(n136), .Y(n140) );
  AOI22XL U244 ( .A0(n27), .A1(n505), .B0(n16), .B1(n504), .Y(n506) );
  NAND2XL U245 ( .A(n6), .B(n37), .Y(n404) );
  OAI2BB1XL U246 ( .A0N(b[1]), .A1N(n43), .B0(n540), .Y(n359) );
  INVXL U247 ( .A(b[0]), .Y(n362) );
  AND2X1 U248 ( .A(n33), .B(b[2]), .Y(n422) );
  XOR3X2 U249 ( .A(n374), .B(n58), .C(n1), .Y(n375) );
  OR2X2 U250 ( .A(n385), .B(n380), .Y(n77) );
  XOR3X2 U251 ( .A(n61), .B(n77), .C(n416), .Y(n377) );
  XOR2X1 U252 ( .A(n559), .B(n3), .Y(n353) );
  XNOR3X2 U253 ( .A(n530), .B(n298), .C(n297), .Y(n299) );
  XOR2X1 U254 ( .A(n339), .B(n290), .Y(n300) );
  XNOR3X2 U255 ( .A(n179), .B(n178), .C(n177), .Y(n192) );
  XOR3X2 U256 ( .A(n81), .B(n374), .C(n416), .Y(n204) );
  XOR2X1 U257 ( .A(n325), .B(n373), .Y(n83) );
  CLKINVX3 U258 ( .A(n152), .Y(n374) );
  XOR2X1 U259 ( .A(n456), .B(n455), .Y(c[12]) );
  XOR2X1 U260 ( .A(n454), .B(n453), .Y(n455) );
  XOR2X1 U261 ( .A(n448), .B(n447), .Y(n456) );
  XOR2X1 U262 ( .A(n450), .B(n449), .Y(n454) );
  XOR2X1 U263 ( .A(n259), .B(n254), .Y(c[6]) );
  XNOR3X2 U264 ( .A(n372), .B(n526), .C(n205), .Y(n259) );
  XOR2X1 U265 ( .A(n84), .B(n1), .Y(n254) );
  XOR2X1 U266 ( .A(n355), .B(n516), .Y(n205) );
  XOR3X2 U267 ( .A(n494), .B(n489), .C(n372), .Y(n497) );
  NOR2X1 U268 ( .A(n381), .B(n400), .Y(n489) );
  XNOR3X2 U269 ( .A(n85), .B(n353), .C(n86), .Y(c[11]) );
  XNOR3X2 U270 ( .A(n431), .B(n352), .C(n351), .Y(n85) );
  AOI22X1 U271 ( .A0(a[0]), .A1(n458), .B0(a[1]), .B1(n457), .Y(n463) );
  OAI21XL U272 ( .A0(a[1]), .A1(n12), .B0(n551), .Y(n458) );
  OAI21XL U273 ( .A0(n102), .A1(n553), .B0(n10), .Y(n457) );
  OAI21XL U274 ( .A0(n108), .A1(n12), .B0(n111), .Y(n518) );
  OAI21XL U275 ( .A0(n107), .A1(n362), .B0(n64), .Y(n517) );
  AOI22X1 U276 ( .A0(n103), .A1(n465), .B0(n25), .B1(n464), .Y(n467) );
  OAI21XL U277 ( .A0(n104), .A1(n12), .B0(n111), .Y(n465) );
  OAI21XL U278 ( .A0(n103), .A1(n362), .B0(n64), .Y(n464) );
  OAI21XL U279 ( .A0(n30), .A1(n12), .B0(n111), .Y(n528) );
  OAI21XL U280 ( .A0(n28), .A1(n362), .B0(n64), .Y(n527) );
  OAI21XL U281 ( .A0(n106), .A1(n12), .B0(n111), .Y(n499) );
  OAI21XL U282 ( .A0(n105), .A1(n362), .B0(n64), .Y(n498) );
  NOR2X1 U283 ( .A(n540), .B(n519), .Y(n520) );
  OAI2BB1X1 U284 ( .A0N(n50), .A1N(n305), .B0(n304), .Y(n306) );
  OAI21XL U285 ( .A0(n9), .A1(n362), .B0(n64), .Y(n421) );
  OAI21XL U286 ( .A0(n33), .A1(n12), .B0(n111), .Y(n538) );
  OAI21XL U287 ( .A0(n30), .A1(n362), .B0(n64), .Y(n537) );
  OAI21XL U288 ( .A0(n27), .A1(n362), .B0(n64), .Y(n504) );
  OAI21XL U289 ( .A0(n104), .A1(n362), .B0(n64), .Y(n490) );
  OAI21XL U290 ( .A0(n37), .A1(n12), .B0(n111), .Y(n420) );
  OAI2BB1X1 U291 ( .A0N(n24), .A1N(n150), .B0(n149), .Y(n151) );
  OAI21XL U292 ( .A0(n148), .A1(n364), .B0(n11), .Y(n149) );
  XOR2X2 U293 ( .A(n175), .B(n174), .Y(n372) );
  XNOR3X2 U294 ( .A(n485), .B(n486), .C(n162), .Y(n175) );
  XNOR3X2 U295 ( .A(n173), .B(n170), .C(n169), .Y(n174) );
  INVX1 U296 ( .A(n100), .Y(n239) );
  NAND2BX1 U297 ( .AN(n14), .B(n43), .Y(n240) );
  INVX1 U298 ( .A(b[11]), .Y(n126) );
  OAI21XL U299 ( .A0(n180), .A1(n302), .B0(n19), .Y(n181) );
  NOR2BX1 U300 ( .AN(n110), .B(n100), .Y(n180) );
  OAI21XL U301 ( .A0(n303), .A1(n302), .B0(n23), .Y(n304) );
  XOR2X1 U302 ( .A(n217), .B(n216), .Y(n219) );
  XNOR3X2 U303 ( .A(n215), .B(n214), .C(n213), .Y(n220) );
  NOR2BX1 U304 ( .AN(n38), .B(n24), .Y(n148) );
  NOR2BX1 U305 ( .AN(n110), .B(n18), .Y(n166) );
  NAND2X1 U306 ( .A(n106), .B(b[11]), .Y(n476) );
  NAND2X1 U307 ( .A(n104), .B(n5), .Y(n522) );
  XOR2X1 U308 ( .A(n314), .B(n311), .Y(n316) );
  NAND2X1 U309 ( .A(n108), .B(n101), .Y(n221) );
  XNOR3X2 U310 ( .A(n355), .B(n426), .C(n87), .Y(n356) );
  XOR2X1 U311 ( .A(n427), .B(n354), .Y(n87) );
  XNOR3X2 U312 ( .A(n501), .B(n202), .C(n195), .Y(n203) );
  XNOR3X2 U313 ( .A(n324), .B(n84), .C(n323), .Y(c[9]) );
  XNOR3X2 U314 ( .A(n316), .B(n315), .C(n559), .Y(n324) );
  XOR3X2 U315 ( .A(n557), .B(n558), .C(n319), .Y(n321) );
  XOR2X1 U316 ( .A(n414), .B(n413), .Y(n415) );
  XOR2X1 U317 ( .A(n410), .B(n409), .Y(n414) );
  XOR2X1 U318 ( .A(n525), .B(n524), .Y(n526) );
  XOR2X1 U319 ( .A(n523), .B(n522), .Y(n524) );
  XOR2X1 U320 ( .A(n521), .B(n520), .Y(n525) );
  XNOR2X1 U321 ( .A(n373), .B(n92), .Y(n376) );
  XNOR2X1 U322 ( .A(n446), .B(n559), .Y(n447) );
  XOR3X2 U323 ( .A(n251), .B(n250), .C(n249), .Y(n252) );
  NAND2X1 U324 ( .A(a[7]), .B(n24), .Y(n249) );
  NAND2X1 U325 ( .A(b[8]), .B(n36), .Y(n250) );
  NAND2X1 U326 ( .A(b[9]), .B(n8), .Y(n251) );
  XOR2X1 U327 ( .A(n546), .B(n545), .Y(n547) );
  XNOR3X2 U328 ( .A(n1), .B(n373), .C(n153), .Y(c[2]) );
  XOR2X1 U329 ( .A(n152), .B(n484), .Y(n153) );
  XOR2X1 U330 ( .A(n467), .B(n466), .Y(n484) );
  NOR2X1 U331 ( .A(n381), .B(n540), .Y(n466) );
  XNOR3X2 U332 ( .A(n461), .B(n145), .C(n144), .Y(n146) );
  XNOR3X2 U333 ( .A(n141), .B(n140), .C(n139), .Y(n147) );
  XOR2X1 U334 ( .A(n406), .B(n405), .Y(n407) );
  XOR2X1 U335 ( .A(n412), .B(n411), .Y(n413) );
  XOR2X1 U336 ( .A(n436), .B(n435), .Y(n437) );
  XOR2X1 U337 ( .A(n479), .B(n478), .Y(n480) );
  XOR2X1 U338 ( .A(n475), .B(n474), .Y(n479) );
  XOR2X1 U339 ( .A(n477), .B(n476), .Y(n478) );
  XNOR3X2 U340 ( .A(n350), .B(n349), .C(n348), .Y(n351) );
  XNOR2X1 U341 ( .A(n347), .B(n346), .Y(n348) );
  XOR3X2 U342 ( .A(n423), .B(n327), .C(n326), .Y(n337) );
  INVX1 U343 ( .A(n105), .Y(n481) );
  OAI2BB1X1 U344 ( .A0N(n23), .A1N(n266), .B0(n265), .Y(n286) );
  OAI21XL U345 ( .A0(n264), .A1(n302), .B0(n21), .Y(n265) );
  NOR2BX1 U346 ( .AN(n110), .B(n99), .Y(n135) );
  XOR3X2 U347 ( .A(n95), .B(n138), .C(n460), .Y(n139) );
  XOR3X2 U348 ( .A(n332), .B(n331), .C(n330), .Y(n333) );
  XOR2X1 U349 ( .A(n262), .B(n261), .Y(n288) );
  XNOR3X2 U350 ( .A(n339), .B(n83), .C(n338), .Y(c[10]) );
  XNOR3X2 U351 ( .A(n335), .B(n334), .C(n333), .Y(n336) );
  INVX1 U352 ( .A(n103), .Y(n380) );
  OAI2BB1X1 U353 ( .A0N(n19), .A1N(n168), .B0(n167), .Y(n169) );
  XOR2X1 U354 ( .A(n542), .B(n541), .Y(n546) );
  NOR2X1 U355 ( .A(n540), .B(n539), .Y(n541) );
  XOR2X1 U356 ( .A(n535), .B(n534), .Y(n536) );
  XOR2X1 U357 ( .A(n445), .B(n444), .Y(n448) );
  XOR2X1 U358 ( .A(n443), .B(n442), .Y(n444) );
  XOR2X1 U359 ( .A(n438), .B(n437), .Y(n445) );
  XOR2X1 U360 ( .A(n441), .B(n440), .Y(n442) );
  NOR2X1 U361 ( .A(n381), .B(n553), .Y(n419) );
  OAI2BB1X1 U362 ( .A0N(n100), .A1N(n182), .B0(n181), .Y(n187) );
  XOR2X1 U363 ( .A(n318), .B(n317), .Y(n319) );
  XOR2X1 U364 ( .A(n513), .B(n512), .Y(c[5]) );
  XOR2X1 U365 ( .A(n511), .B(n510), .Y(n513) );
  XOR2X1 U366 ( .A(n509), .B(n508), .Y(n510) );
  XOR2X1 U367 ( .A(n493), .B(n492), .Y(n494) );
  NOR2X1 U368 ( .A(n380), .B(n540), .Y(n492) );
  AOI22X1 U369 ( .A0(n104), .A1(n491), .B0(n26), .B1(n490), .Y(n493) );
  OAI21XL U370 ( .A0(n105), .A1(n12), .B0(n111), .Y(n491) );
  XOR2X1 U371 ( .A(n425), .B(n424), .Y(n335) );
  XNOR2X1 U372 ( .A(n462), .B(n459), .Y(n144) );
  OAI21XL U373 ( .A0(n38), .A1(n552), .B0(n111), .Y(n430) );
  OAI21XL U374 ( .A0(n37), .A1(n362), .B0(n10), .Y(n429) );
  OAI21XL U375 ( .A0(n9), .A1(n12), .B0(n551), .Y(n555) );
  OAI21XL U376 ( .A0(n33), .A1(n553), .B0(n10), .Y(n554) );
  XOR2X1 U377 ( .A(n487), .B(n488), .Y(n162) );
  NOR2X1 U378 ( .A(n540), .B(n378), .Y(n529) );
  XOR2X1 U379 ( .A(n452), .B(n451), .Y(n453) );
  XOR2X1 U380 ( .A(n434), .B(n433), .Y(n352) );
  XOR2X1 U381 ( .A(n544), .B(n543), .Y(n545) );
  XOR2X1 U382 ( .A(n515), .B(n514), .Y(n516) );
  XNOR3X2 U383 ( .A(n532), .B(n296), .C(n295), .Y(n297) );
  INVX1 U384 ( .A(n102), .Y(n381) );
  XOR2X1 U385 ( .A(n194), .B(n500), .Y(n195) );
  NAND2X1 U386 ( .A(n102), .B(n5), .Y(n194) );
  NOR2X1 U387 ( .A(n540), .B(n550), .Y(n500) );
  INVX1 U388 ( .A(n104), .Y(n550) );
  MXI2X1 U389 ( .A(n361), .B(n358), .S0(b[1]), .Y(n360) );
  NAND2XL U390 ( .A(n98), .B(n134), .Y(n137) );
  OAI21XL U391 ( .A0(n135), .A1(n302), .B0(b[2]), .Y(n136) );
  BUFX3 U392 ( .A(a[6]), .Y(n108) );
  BUFX3 U393 ( .A(a[2]), .Y(n104) );
  XOR2X1 U394 ( .A(n96), .B(n97), .Y(n315) );
  BUFX3 U395 ( .A(a[3]), .Y(n105) );
  BUFX3 U396 ( .A(a[5]), .Y(n107) );
  BUFX3 U397 ( .A(a[4]), .Y(n106) );
  BUFX3 U398 ( .A(a[1]), .Y(n103) );
  INVX1 U399 ( .A(b[0]), .Y(n553) );
  INVX1 U400 ( .A(b[1]), .Y(n552) );
  BUFX3 U401 ( .A(b[12]), .Y(n101) );
  BUFX3 U402 ( .A(n551), .Y(n111) );
  XOR2X1 U403 ( .A(n507), .B(n506), .Y(n511) );
  OAI21XL U404 ( .A0(n16), .A1(n12), .B0(n111), .Y(n505) );
  XOR2X1 U405 ( .A(n404), .B(n403), .Y(n408) );
  OAI21X1 U406 ( .A0(n360), .A1(n364), .B0(n359), .Y(n403) );
  XOR2X1 U407 ( .A(n366), .B(n439), .Y(n443) );
  AOI2BB2X1 U408 ( .B0(b[1]), .B1(n364), .A0N(n357), .A1N(n362), .Y(n365) );
  BUFX3 U409 ( .A(a[0]), .Y(n102) );
  XOR2X1 U410 ( .A(n204), .B(n463), .Y(c[1]) );
  NAND2X1 U411 ( .A(n26), .B(b[2]), .Y(n507) );
  NAND2X1 U412 ( .A(b[2]), .B(n37), .Y(n439) );
  NAND2BXL U413 ( .AN(b[2]), .B(n109), .Y(n134) );
  NAND2BX4 U414 ( .AN(n110), .B(n109), .Y(n368) );
  AND2X4 U415 ( .A(n8), .B(n18), .Y(n138) );
endmodule


module feedback_ckt_15 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  mux_13_18 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX1 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
endmodule


module feedback_ckt_14 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;
  wire   n1;
  wire   [12:0] out;

  DFFRHQX4 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  mux_13_17 mux ( .a({Qout[12], n1, Qout[10:0]}), .b(Din), .sel(start), .out(
        out) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX4 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  BUFX3 U3 ( .A(Qout[11]), .Y(n1) );
endmodule


module feedback_ckt_13 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  mux_13_16 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX1 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
endmodule


module feedback_ckt_12 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  DFFRHQX4 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX4 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  mux_13_15 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
endmodule


module feedback_ckt_11 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  mux_13_13 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX1 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX2 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
endmodule


module feedback_ckt_10 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  DFFRHQX4 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX4 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  mux_13_12 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
endmodule


module feedback_ckt_9 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  mux_13_11 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX1 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
endmodule


module feedback_ckt_8 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  DFFRHQX4 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  mux_13_10 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX4 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
endmodule


module feedback_ckt_7 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;
  wire   n2;
  wire   [12:0] out;

  mux_13_8 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(n2) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX1 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX2 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  BUFX3 U3 ( .A(n2), .Y(Qout[4]) );
endmodule


module feedback_ckt_6 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  mux_13_7 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX4 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  DFFRHQX2 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
endmodule


module feedback_ckt_5 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  mux_13_6 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX1 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
endmodule


module feedback_ckt_4 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  DFFRHQX4 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  mux_13_5 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX4 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
endmodule


module feedback_ckt_3 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  mux_13_3 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX1 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
endmodule


module feedback_ckt_2 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  DFFRHQX4 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  mux_13_2 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX4 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
endmodule


module feedback_ckt_1 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  mux_13_1 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX1 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
endmodule


module feedback_ckt_0 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  DFFRHQX4 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX4 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  mux_13_0 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
endmodule


module degree_computation_2 ( deg_Ri, deg_Qi, stop_i, d1out, start, deg_Ro, 
        deg_Qo, stop_o, sw, clk, reset );
  input [4:0] deg_Ri;
  input [4:0] deg_Qi;
  input [12:0] d1out;
  output [4:0] deg_Ro;
  output [4:0] deg_Qo;
  input stop_i, start, clk, reset;
  output stop_o, sw;
  wire   out, sw_reg, stop2_signal, n1, n7, n8, n9, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [4:0] DQ1;
  wire   [4:0] DR1;
  wire   [4:0] rmux_signal;
  wire   [4:0] qmux_signal;
  wire   [4:0] DR2;
  wire   [4:0] addr_signal;
  wire   [4:0] DQ2;
  wire   [4:0] addq_signal;
  wire   [4:0] mr_signal;
  wire   [4:0] mq_signal;
  wire   [4:0] r2mux_signal;
  wire   [4:0] q2mux_signal;
  wire   [12:0] dmux_signal;

  mux_5_17 mdeg1 ( .a(DQ1), .b(DR1), .sel(n9), .out(rmux_signal) );
  mux_5_16 mdeg2 ( .a(DR1), .b(DQ1), .sel(sw_reg), .out(qmux_signal) );
  mux_5_15 mdeg3 ( .a(DR2), .b(addr_signal), .sel(n8), .out(mr_signal) );
  mux_5_14 mdeg4 ( .a(addq_signal), .b(DQ2), .sel(n7), .out(mq_signal) );
  mux_5_13 mdeg5 ( .a(DR2), .b(mr_signal), .sel(n11), .out(r2mux_signal) );
  mux_5_12 mdeg6 ( .a(DQ2), .b(mq_signal), .sel(n11), .out(q2mux_signal) );
  mux_13_14 mdeg7 ( .a(d1out), .b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .sel(stop2_signal), .out(
        dmux_signal) );
  degree_computation_2_DW01_dec_0 sub_41 ( .A(DQ2), .SUM(addq_signal) );
  degree_computation_2_DW01_dec_1 sub_40 ( .A(DR2), .SUM(addr_signal) );
  DFFRHQX1 \DQ3_reg[2]  ( .D(q2mux_signal[2]), .CK(clk), .RN(reset), .Q(
        deg_Qo[2]) );
  DFFRHQX1 \DQ3_reg[3]  ( .D(q2mux_signal[3]), .CK(clk), .RN(reset), .Q(
        deg_Qo[3]) );
  DFFRHQX1 \DQ3_reg[4]  ( .D(q2mux_signal[4]), .CK(clk), .RN(reset), .Q(
        deg_Qo[4]) );
  DFFRHQX1 \DR3_reg[1]  ( .D(r2mux_signal[1]), .CK(clk), .RN(reset), .Q(
        deg_Ro[1]) );
  DFFRHQX1 \DR3_reg[0]  ( .D(r2mux_signal[0]), .CK(clk), .RN(reset), .Q(
        deg_Ro[0]) );
  DFFRHQX1 \DQ3_reg[0]  ( .D(q2mux_signal[0]), .CK(clk), .RN(reset), .Q(
        deg_Qo[0]) );
  DFFRHQX1 \DR3_reg[3]  ( .D(r2mux_signal[3]), .CK(clk), .RN(reset), .Q(
        deg_Ro[3]) );
  DFFRHQX1 \DR3_reg[4]  ( .D(r2mux_signal[4]), .CK(clk), .RN(reset), .Q(
        deg_Ro[4]) );
  DFFRHQX1 \DQ3_reg[1]  ( .D(q2mux_signal[1]), .CK(clk), .RN(reset), .Q(
        deg_Qo[1]) );
  DFFRHQX1 \DR3_reg[2]  ( .D(r2mux_signal[2]), .CK(clk), .RN(reset), .Q(
        deg_Ro[2]) );
  DFFRHQX1 \DQ1_reg[3]  ( .D(deg_Qi[3]), .CK(clk), .RN(reset), .Q(DQ1[3]) );
  DFFRHQX1 \DQ1_reg[2]  ( .D(deg_Qi[2]), .CK(clk), .RN(reset), .Q(DQ1[2]) );
  DFFRHQX1 \DQ1_reg[1]  ( .D(deg_Qi[1]), .CK(clk), .RN(reset), .Q(DQ1[1]) );
  DFFRHQX1 \DQ1_reg[0]  ( .D(deg_Qi[0]), .CK(clk), .RN(reset), .Q(DQ1[0]) );
  DFFRHQX1 \DR1_reg[3]  ( .D(deg_Ri[3]), .CK(clk), .RN(reset), .Q(DR1[3]) );
  DFFRHQX1 \DR1_reg[2]  ( .D(deg_Ri[2]), .CK(clk), .RN(reset), .Q(DR1[2]) );
  DFFRHQX1 \DR1_reg[1]  ( .D(deg_Ri[1]), .CK(clk), .RN(reset), .Q(DR1[1]) );
  DFFRHQX1 \DR1_reg[0]  ( .D(deg_Ri[0]), .CK(clk), .RN(reset), .Q(DR1[0]) );
  DFFRHQX1 \DQ1_reg[4]  ( .D(deg_Qi[4]), .CK(clk), .RN(reset), .Q(DQ1[4]) );
  DFFRHQX1 \DR1_reg[4]  ( .D(deg_Ri[4]), .CK(clk), .RN(reset), .Q(DR1[4]) );
  DFFRHQX1 \DQ2_reg[4]  ( .D(qmux_signal[4]), .CK(clk), .RN(reset), .Q(DQ2[4])
         );
  DFFRHQX1 \DR2_reg[4]  ( .D(rmux_signal[4]), .CK(clk), .RN(reset), .Q(DR2[4])
         );
  DFFRHQX1 sw_reg_reg ( .D(out), .CK(clk), .RN(reset), .Q(sw_reg) );
  DFFRHQX1 shift_reg_reg ( .D(out), .CK(clk), .RN(reset), .Q(sw) );
  DFFRHQX1 \DQ2_reg[2]  ( .D(qmux_signal[2]), .CK(clk), .RN(reset), .Q(DQ2[2])
         );
  DFFRHQX1 \DR2_reg[2]  ( .D(rmux_signal[2]), .CK(clk), .RN(reset), .Q(DR2[2])
         );
  DFFRHQX1 \DQ2_reg[1]  ( .D(qmux_signal[1]), .CK(clk), .RN(reset), .Q(DQ2[1])
         );
  DFFRHQX1 \DR2_reg[1]  ( .D(rmux_signal[1]), .CK(clk), .RN(reset), .Q(DR2[1])
         );
  DFFRHQX1 \DQ2_reg[3]  ( .D(qmux_signal[3]), .CK(clk), .RN(reset), .Q(DQ2[3])
         );
  DFFRHQX1 \DR2_reg[3]  ( .D(rmux_signal[3]), .CK(clk), .RN(reset), .Q(DR2[3])
         );
  DFFRHQX1 \DQ2_reg[0]  ( .D(qmux_signal[0]), .CK(clk), .RN(reset), .Q(DQ2[0])
         );
  DFFRHQX1 \DR2_reg[0]  ( .D(rmux_signal[0]), .CK(clk), .RN(reset), .Q(DR2[0])
         );
  DFFSX1 start_reg_reg ( .D(start), .CK(clk), .SN(reset), .Q(stop2_signal) );
  NAND4X1 U3 ( .A(n26), .B(n25), .C(n24), .D(n23), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n7) );
  INVX1 U5 ( .A(n1), .Y(n8) );
  BUFX3 U6 ( .A(sw_reg), .Y(n9) );
  INVX1 U7 ( .A(n12), .Y(n11) );
  INVX1 U8 ( .A(stop_i), .Y(n12) );
  NOR3X1 U9 ( .A(dmux_signal[0]), .B(dmux_signal[11]), .C(dmux_signal[10]), 
        .Y(n26) );
  NOR3X1 U10 ( .A(dmux_signal[12]), .B(dmux_signal[2]), .C(dmux_signal[1]), 
        .Y(n25) );
  NOR3X1 U11 ( .A(dmux_signal[3]), .B(dmux_signal[5]), .C(dmux_signal[4]), .Y(
        n24) );
  NOR4X1 U12 ( .A(dmux_signal[9]), .B(dmux_signal[8]), .C(dmux_signal[7]), .D(
        dmux_signal[6]), .Y(n23) );
  AND2X2 U13 ( .A(stop2_signal), .B(n27), .Y(stop_o) );
  OAI22X1 U14 ( .A0(mr_signal[4]), .A1(mr_signal[3]), .B0(mq_signal[4]), .B1(
        mq_signal[3]), .Y(n27) );
  INVX1 U15 ( .A(deg_Qi[4]), .Y(n22) );
  INVX1 U16 ( .A(deg_Ri[1]), .Y(n15) );
  AOI2BB1X1 U17 ( .A0N(n15), .A1N(deg_Qi[1]), .B0(deg_Ri[0]), .Y(n14) );
  INVX1 U18 ( .A(deg_Qi[2]), .Y(n17) );
  INVX1 U19 ( .A(deg_Qi[3]), .Y(n13) );
  AND2X1 U20 ( .A(deg_Ri[3]), .B(n13), .Y(n16) );
  OAI32X1 U21 ( .A0(n17), .A1(deg_Ri[2]), .A2(n16), .B0(deg_Ri[3]), .B1(n13), 
        .Y(n18) );
  AOI221X1 U22 ( .A0(deg_Qi[1]), .A1(n15), .B0(n14), .B1(deg_Qi[0]), .C0(n18), 
        .Y(n21) );
  AOI21X1 U23 ( .A0(deg_Ri[2]), .A1(n17), .B0(n16), .Y(n19) );
  OAI2BB2X1 U24 ( .B0(n19), .B1(n18), .A0N(n22), .A1N(deg_Ri[4]), .Y(n20) );
  OAI22X1 U25 ( .A0(deg_Ri[4]), .A1(n22), .B0(n21), .B1(n20), .Y(out) );
endmodule


module degree_computation_1 ( deg_Ri, deg_Qi, stop_i, d1out, start, deg_Ro, 
        deg_Qo, stop_o, sw, clk, reset );
  input [4:0] deg_Ri;
  input [4:0] deg_Qi;
  input [12:0] d1out;
  output [4:0] deg_Ro;
  output [4:0] deg_Qo;
  input stop_i, start, clk, reset;
  output stop_o, sw;
  wire   out, sw_reg, stop2_signal, n1, n7, n8, n9, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [4:0] DQ1;
  wire   [4:0] DR1;
  wire   [4:0] rmux_signal;
  wire   [4:0] qmux_signal;
  wire   [4:0] DR2;
  wire   [4:0] addr_signal;
  wire   [4:0] DQ2;
  wire   [4:0] addq_signal;
  wire   [4:0] mr_signal;
  wire   [4:0] mq_signal;
  wire   [4:0] r2mux_signal;
  wire   [4:0] q2mux_signal;
  wire   [12:0] dmux_signal;

  mux_5_11 mdeg1 ( .a(DQ1), .b(DR1), .sel(n9), .out(rmux_signal) );
  mux_5_10 mdeg2 ( .a(DR1), .b(DQ1), .sel(sw_reg), .out(qmux_signal) );
  mux_5_9 mdeg3 ( .a(DR2), .b(addr_signal), .sel(n8), .out(mr_signal) );
  mux_5_8 mdeg4 ( .a(addq_signal), .b(DQ2), .sel(n7), .out(mq_signal) );
  mux_5_7 mdeg5 ( .a(DR2), .b(mr_signal), .sel(n11), .out(r2mux_signal) );
  mux_5_6 mdeg6 ( .a(DQ2), .b(mq_signal), .sel(n11), .out(q2mux_signal) );
  mux_13_9 mdeg7 ( .a(d1out), .b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .sel(stop2_signal), .out(
        dmux_signal) );
  degree_computation_1_DW01_dec_0 sub_41 ( .A(DQ2), .SUM(addq_signal) );
  degree_computation_1_DW01_dec_1 sub_40 ( .A(DR2), .SUM(addr_signal) );
  DFFRHQX1 \DQ3_reg[2]  ( .D(q2mux_signal[2]), .CK(clk), .RN(reset), .Q(
        deg_Qo[2]) );
  DFFRHQX1 \DQ3_reg[3]  ( .D(q2mux_signal[3]), .CK(clk), .RN(reset), .Q(
        deg_Qo[3]) );
  DFFRHQX1 \DQ3_reg[4]  ( .D(q2mux_signal[4]), .CK(clk), .RN(reset), .Q(
        deg_Qo[4]) );
  DFFRHQX1 \DR3_reg[1]  ( .D(r2mux_signal[1]), .CK(clk), .RN(reset), .Q(
        deg_Ro[1]) );
  DFFRHQX1 \DR3_reg[0]  ( .D(r2mux_signal[0]), .CK(clk), .RN(reset), .Q(
        deg_Ro[0]) );
  DFFRHQX1 \DQ3_reg[0]  ( .D(q2mux_signal[0]), .CK(clk), .RN(reset), .Q(
        deg_Qo[0]) );
  DFFRHQX1 \DR3_reg[3]  ( .D(r2mux_signal[3]), .CK(clk), .RN(reset), .Q(
        deg_Ro[3]) );
  DFFRHQX1 \DR3_reg[4]  ( .D(r2mux_signal[4]), .CK(clk), .RN(reset), .Q(
        deg_Ro[4]) );
  DFFRHQX1 \DQ3_reg[1]  ( .D(q2mux_signal[1]), .CK(clk), .RN(reset), .Q(
        deg_Qo[1]) );
  DFFRHQX1 \DR3_reg[2]  ( .D(r2mux_signal[2]), .CK(clk), .RN(reset), .Q(
        deg_Ro[2]) );
  DFFRHQX1 \DQ1_reg[3]  ( .D(deg_Qi[3]), .CK(clk), .RN(reset), .Q(DQ1[3]) );
  DFFRHQX1 \DQ1_reg[2]  ( .D(deg_Qi[2]), .CK(clk), .RN(reset), .Q(DQ1[2]) );
  DFFRHQX1 \DQ1_reg[1]  ( .D(deg_Qi[1]), .CK(clk), .RN(reset), .Q(DQ1[1]) );
  DFFRHQX1 \DQ1_reg[0]  ( .D(deg_Qi[0]), .CK(clk), .RN(reset), .Q(DQ1[0]) );
  DFFRHQX1 \DR1_reg[3]  ( .D(deg_Ri[3]), .CK(clk), .RN(reset), .Q(DR1[3]) );
  DFFRHQX1 \DR1_reg[2]  ( .D(deg_Ri[2]), .CK(clk), .RN(reset), .Q(DR1[2]) );
  DFFRHQX1 \DR1_reg[1]  ( .D(deg_Ri[1]), .CK(clk), .RN(reset), .Q(DR1[1]) );
  DFFRHQX1 \DR1_reg[0]  ( .D(deg_Ri[0]), .CK(clk), .RN(reset), .Q(DR1[0]) );
  DFFRHQX1 \DQ1_reg[4]  ( .D(deg_Qi[4]), .CK(clk), .RN(reset), .Q(DQ1[4]) );
  DFFRHQX1 \DR1_reg[4]  ( .D(deg_Ri[4]), .CK(clk), .RN(reset), .Q(DR1[4]) );
  DFFRHQX1 \DQ2_reg[4]  ( .D(qmux_signal[4]), .CK(clk), .RN(reset), .Q(DQ2[4])
         );
  DFFRHQX1 \DR2_reg[4]  ( .D(rmux_signal[4]), .CK(clk), .RN(reset), .Q(DR2[4])
         );
  DFFRHQX1 sw_reg_reg ( .D(out), .CK(clk), .RN(reset), .Q(sw_reg) );
  DFFRHQX1 shift_reg_reg ( .D(out), .CK(clk), .RN(reset), .Q(sw) );
  DFFRHQX1 \DQ2_reg[2]  ( .D(qmux_signal[2]), .CK(clk), .RN(reset), .Q(DQ2[2])
         );
  DFFRHQX1 \DR2_reg[2]  ( .D(rmux_signal[2]), .CK(clk), .RN(reset), .Q(DR2[2])
         );
  DFFRHQX1 \DQ2_reg[1]  ( .D(qmux_signal[1]), .CK(clk), .RN(reset), .Q(DQ2[1])
         );
  DFFRHQX1 \DR2_reg[1]  ( .D(rmux_signal[1]), .CK(clk), .RN(reset), .Q(DR2[1])
         );
  DFFRHQX1 \DQ2_reg[3]  ( .D(qmux_signal[3]), .CK(clk), .RN(reset), .Q(DQ2[3])
         );
  DFFRHQX1 \DR2_reg[3]  ( .D(rmux_signal[3]), .CK(clk), .RN(reset), .Q(DR2[3])
         );
  DFFRHQX1 \DQ2_reg[0]  ( .D(qmux_signal[0]), .CK(clk), .RN(reset), .Q(DQ2[0])
         );
  DFFRHQX1 \DR2_reg[0]  ( .D(rmux_signal[0]), .CK(clk), .RN(reset), .Q(DR2[0])
         );
  DFFSX1 start_reg_reg ( .D(start), .CK(clk), .SN(reset), .Q(stop2_signal) );
  NAND4X1 U3 ( .A(n26), .B(n25), .C(n24), .D(n23), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n7) );
  INVX1 U5 ( .A(n1), .Y(n8) );
  BUFX3 U6 ( .A(sw_reg), .Y(n9) );
  INVX1 U7 ( .A(n12), .Y(n11) );
  INVX1 U8 ( .A(stop_i), .Y(n12) );
  NOR3X1 U9 ( .A(dmux_signal[0]), .B(dmux_signal[11]), .C(dmux_signal[10]), 
        .Y(n26) );
  NOR3X1 U10 ( .A(dmux_signal[12]), .B(dmux_signal[2]), .C(dmux_signal[1]), 
        .Y(n25) );
  NOR3X1 U11 ( .A(dmux_signal[3]), .B(dmux_signal[5]), .C(dmux_signal[4]), .Y(
        n24) );
  NOR4X1 U12 ( .A(dmux_signal[9]), .B(dmux_signal[8]), .C(dmux_signal[7]), .D(
        dmux_signal[6]), .Y(n23) );
  AND2X2 U13 ( .A(stop2_signal), .B(n27), .Y(stop_o) );
  OAI22X1 U14 ( .A0(mr_signal[4]), .A1(mr_signal[3]), .B0(mq_signal[4]), .B1(
        mq_signal[3]), .Y(n27) );
  INVX1 U15 ( .A(deg_Qi[4]), .Y(n22) );
  INVX1 U16 ( .A(deg_Ri[1]), .Y(n15) );
  AOI2BB1X1 U17 ( .A0N(n15), .A1N(deg_Qi[1]), .B0(deg_Ri[0]), .Y(n14) );
  INVX1 U18 ( .A(deg_Qi[2]), .Y(n17) );
  INVX1 U19 ( .A(deg_Qi[3]), .Y(n13) );
  AND2X1 U20 ( .A(deg_Ri[3]), .B(n13), .Y(n16) );
  OAI32X1 U21 ( .A0(n17), .A1(deg_Ri[2]), .A2(n16), .B0(deg_Ri[3]), .B1(n13), 
        .Y(n18) );
  AOI221X1 U22 ( .A0(deg_Qi[1]), .A1(n15), .B0(n14), .B1(deg_Qi[0]), .C0(n18), 
        .Y(n21) );
  AOI21X1 U23 ( .A0(deg_Ri[2]), .A1(n17), .B0(n16), .Y(n19) );
  OAI2BB2X1 U24 ( .B0(n19), .B1(n18), .A0N(n22), .A1N(deg_Ri[4]), .Y(n20) );
  OAI22X1 U25 ( .A0(deg_Ri[4]), .A1(n22), .B0(n21), .B1(n20), .Y(out) );
endmodule


module degree_computation_0 ( deg_Ri, deg_Qi, stop_i, d1out, start, deg_Ro, 
        deg_Qo, stop_o, sw, clk, reset );
  input [4:0] deg_Ri;
  input [4:0] deg_Qi;
  input [12:0] d1out;
  output [4:0] deg_Ro;
  output [4:0] deg_Qo;
  input stop_i, start, clk, reset;
  output stop_o, sw;
  wire   out, sw_reg, stop2_signal, n1, n7, n8, n9, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;
  wire   [4:0] DQ1;
  wire   [4:0] DR1;
  wire   [4:0] rmux_signal;
  wire   [4:0] qmux_signal;
  wire   [4:0] DR2;
  wire   [4:0] addr_signal;
  wire   [4:0] DQ2;
  wire   [4:0] addq_signal;
  wire   [4:0] mr_signal;
  wire   [4:0] mq_signal;
  wire   [4:0] r2mux_signal;
  wire   [4:0] q2mux_signal;
  wire   [12:0] dmux_signal;

  mux_5_5 mdeg1 ( .a(DQ1), .b(DR1), .sel(n9), .out(rmux_signal) );
  mux_5_4 mdeg2 ( .a(DR1), .b(DQ1), .sel(sw_reg), .out(qmux_signal) );
  mux_5_3 mdeg3 ( .a(DR2), .b(addr_signal), .sel(n8), .out(mr_signal) );
  mux_5_2 mdeg4 ( .a(addq_signal), .b(DQ2), .sel(n7), .out(mq_signal) );
  mux_5_1 mdeg5 ( .a(DR2), .b(mr_signal), .sel(n11), .out(r2mux_signal) );
  mux_5_0 mdeg6 ( .a(DQ2), .b(mq_signal), .sel(n11), .out(q2mux_signal) );
  mux_13_4 mdeg7 ( .a(d1out), .b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .sel(stop2_signal), .out(
        dmux_signal) );
  degree_computation_0_DW01_dec_0 sub_41 ( .A(DQ2), .SUM(addq_signal) );
  degree_computation_0_DW01_dec_1 sub_40 ( .A(DR2), .SUM(addr_signal) );
  DFFRHQX1 \DQ3_reg[0]  ( .D(q2mux_signal[0]), .CK(clk), .RN(reset), .Q(
        deg_Qo[0]) );
  DFFRHQX1 \DQ3_reg[1]  ( .D(q2mux_signal[1]), .CK(clk), .RN(reset), .Q(
        deg_Qo[1]) );
  DFFRHQX1 \DQ3_reg[2]  ( .D(q2mux_signal[2]), .CK(clk), .RN(reset), .Q(
        deg_Qo[2]) );
  DFFRHQX1 \DQ3_reg[3]  ( .D(q2mux_signal[3]), .CK(clk), .RN(reset), .Q(
        deg_Qo[3]) );
  DFFRHQX1 \DQ3_reg[4]  ( .D(q2mux_signal[4]), .CK(clk), .RN(reset), .Q(
        deg_Qo[4]) );
  DFFRHQX1 \DR3_reg[4]  ( .D(r2mux_signal[4]), .CK(clk), .RN(reset), .Q(
        deg_Ro[4]) );
  DFFRHQX1 \DR3_reg[3]  ( .D(r2mux_signal[3]), .CK(clk), .RN(reset), .Q(
        deg_Ro[3]) );
  DFFRHQX1 \DR3_reg[2]  ( .D(r2mux_signal[2]), .CK(clk), .RN(reset), .Q(
        deg_Ro[2]) );
  DFFRHQX1 \DR3_reg[1]  ( .D(r2mux_signal[1]), .CK(clk), .RN(reset), .Q(
        deg_Ro[1]) );
  DFFRHQX1 \DR3_reg[0]  ( .D(r2mux_signal[0]), .CK(clk), .RN(reset), .Q(
        deg_Ro[0]) );
  DFFRHQX1 \DQ1_reg[3]  ( .D(deg_Qi[3]), .CK(clk), .RN(reset), .Q(DQ1[3]) );
  DFFRHQX1 \DQ1_reg[2]  ( .D(deg_Qi[2]), .CK(clk), .RN(reset), .Q(DQ1[2]) );
  DFFRHQX1 \DQ1_reg[1]  ( .D(deg_Qi[1]), .CK(clk), .RN(reset), .Q(DQ1[1]) );
  DFFRHQX1 \DQ1_reg[0]  ( .D(deg_Qi[0]), .CK(clk), .RN(reset), .Q(DQ1[0]) );
  DFFRHQX1 \DR1_reg[3]  ( .D(deg_Ri[3]), .CK(clk), .RN(reset), .Q(DR1[3]) );
  DFFRHQX1 \DR1_reg[2]  ( .D(deg_Ri[2]), .CK(clk), .RN(reset), .Q(DR1[2]) );
  DFFRHQX1 \DR1_reg[1]  ( .D(deg_Ri[1]), .CK(clk), .RN(reset), .Q(DR1[1]) );
  DFFRHQX1 \DR1_reg[0]  ( .D(deg_Ri[0]), .CK(clk), .RN(reset), .Q(DR1[0]) );
  DFFRHQX1 \DQ1_reg[4]  ( .D(deg_Qi[4]), .CK(clk), .RN(reset), .Q(DQ1[4]) );
  DFFRHQX1 \DR1_reg[4]  ( .D(deg_Ri[4]), .CK(clk), .RN(reset), .Q(DR1[4]) );
  DFFRHQX1 sw_reg_reg ( .D(out), .CK(clk), .RN(reset), .Q(sw_reg) );
  DFFRHQX1 shift_reg_reg ( .D(out), .CK(clk), .RN(reset), .Q(sw) );
  DFFRHQX1 \DQ2_reg[2]  ( .D(qmux_signal[2]), .CK(clk), .RN(reset), .Q(DQ2[2])
         );
  DFFRHQX1 \DR2_reg[2]  ( .D(rmux_signal[2]), .CK(clk), .RN(reset), .Q(DR2[2])
         );
  DFFRHQX1 \DQ2_reg[4]  ( .D(qmux_signal[4]), .CK(clk), .RN(reset), .Q(DQ2[4])
         );
  DFFRHQX1 \DR2_reg[4]  ( .D(rmux_signal[4]), .CK(clk), .RN(reset), .Q(DR2[4])
         );
  DFFRHQX1 \DQ2_reg[1]  ( .D(qmux_signal[1]), .CK(clk), .RN(reset), .Q(DQ2[1])
         );
  DFFRHQX1 \DR2_reg[1]  ( .D(rmux_signal[1]), .CK(clk), .RN(reset), .Q(DR2[1])
         );
  DFFRHQX1 \DQ2_reg[3]  ( .D(qmux_signal[3]), .CK(clk), .RN(reset), .Q(DQ2[3])
         );
  DFFRHQX1 \DR2_reg[3]  ( .D(rmux_signal[3]), .CK(clk), .RN(reset), .Q(DR2[3])
         );
  DFFRHQX1 \DQ2_reg[0]  ( .D(qmux_signal[0]), .CK(clk), .RN(reset), .Q(DQ2[0])
         );
  DFFRHQX1 \DR2_reg[0]  ( .D(rmux_signal[0]), .CK(clk), .RN(reset), .Q(DR2[0])
         );
  DFFSX1 start_reg_reg ( .D(start), .CK(clk), .SN(reset), .Q(stop2_signal) );
  NAND4X1 U3 ( .A(n26), .B(n25), .C(n24), .D(n23), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n7) );
  INVX1 U5 ( .A(n1), .Y(n8) );
  BUFX3 U6 ( .A(sw_reg), .Y(n9) );
  INVX1 U7 ( .A(n12), .Y(n11) );
  INVX1 U8 ( .A(stop_i), .Y(n12) );
  NOR3X1 U9 ( .A(dmux_signal[0]), .B(dmux_signal[11]), .C(dmux_signal[10]), 
        .Y(n26) );
  NOR3X1 U10 ( .A(dmux_signal[12]), .B(dmux_signal[2]), .C(dmux_signal[1]), 
        .Y(n25) );
  NOR3X1 U11 ( .A(dmux_signal[3]), .B(dmux_signal[5]), .C(dmux_signal[4]), .Y(
        n24) );
  NOR4X1 U12 ( .A(dmux_signal[9]), .B(dmux_signal[8]), .C(dmux_signal[7]), .D(
        dmux_signal[6]), .Y(n23) );
  AND2X2 U13 ( .A(stop2_signal), .B(n27), .Y(stop_o) );
  OAI22X1 U14 ( .A0(mr_signal[4]), .A1(mr_signal[3]), .B0(mq_signal[4]), .B1(
        mq_signal[3]), .Y(n27) );
  INVX1 U15 ( .A(deg_Qi[4]), .Y(n22) );
  INVX1 U16 ( .A(deg_Ri[1]), .Y(n15) );
  AOI2BB1X1 U17 ( .A0N(n15), .A1N(deg_Qi[1]), .B0(deg_Ri[0]), .Y(n14) );
  INVX1 U18 ( .A(deg_Qi[2]), .Y(n17) );
  INVX1 U19 ( .A(deg_Qi[3]), .Y(n13) );
  AND2X1 U20 ( .A(deg_Ri[3]), .B(n13), .Y(n16) );
  OAI32X1 U21 ( .A0(n17), .A1(deg_Ri[2]), .A2(n16), .B0(deg_Ri[3]), .B1(n13), 
        .Y(n18) );
  AOI221X1 U22 ( .A0(deg_Qi[1]), .A1(n15), .B0(n14), .B1(deg_Qi[0]), .C0(n18), 
        .Y(n21) );
  AOI21X1 U23 ( .A0(deg_Ri[2]), .A1(n17), .B0(n16), .Y(n19) );
  OAI2BB2X1 U24 ( .B0(n19), .B1(n18), .A0N(n22), .A1N(deg_Ri[4]), .Y(n20) );
  OAI22X1 U25 ( .A0(deg_Ri[4]), .A1(n22), .B0(n21), .B1(n20), .Y(out) );
endmodule


module euclidean_cell_2 ( deg_Ri, deg_Qi, stop_i, Rin, Qin, Lin, Uin, start, 
        start_cnt, deg_Ro, deg_Qo, stop_o, Rout, Qout, Lout, Uout, st_out, clk, 
        reset );
  input [4:0] deg_Ri;
  input [4:0] deg_Qi;
  input [12:0] Rin;
  input [12:0] Qin;
  input [12:0] Lin;
  input [12:0] Uin;
  output [4:0] deg_Ro;
  output [4:0] deg_Qo;
  output [12:0] Rout;
  output [12:0] Qout;
  output [12:0] Lout;
  output [12:0] Uout;
  input stop_i, start, start_cnt, clk, reset;
  output stop_o, st_out;
  wire   sw, S2, n2, n57, n58, n61, n62, n63, n64, n65, n122, n123, n124, n126,
         n127, n128, n129, n130, n134, n136, n193, n194, n195, n197, n198,
         n199, n200, n201, n258, n259, n260, n262, n263, n264, n265, n266,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519;
  wire   [12:0] d1out;
  wire   [12:0] Q1;
  wire   [12:0] R1;
  wire   [12:0] r_mux;
  wire   [12:0] q_mux;
  wire   [12:0] U1;
  wire   [12:0] L1;
  wire   [12:0] l_mux;
  wire   [12:0] u_mux;
  wire   [12:0] d2out;
  wire   [12:0] d3out;
  wire   [12:0] d4out;
  wire   [12:0] R2;
  wire   [12:0] m1out;
  wire   [12:0] Q2;
  wire   [12:0] m2out;
  wire   [12:0] L2;
  wire   [12:0] m3out;
  wire   [12:0] U2;
  wire   [12:0] m4out;
  wire   [12:0] add1out;
  wire   [12:0] add2out;
  wire   [12:0] Q3;
  wire   [12:0] U3;

  DFFRHQX4 \R2_reg[12]  ( .D(n331), .CK(clk), .RN(reset), .Q(R2[12]) );
  DFFRHQX4 \L2_reg[12]  ( .D(n388), .CK(clk), .RN(reset), .Q(L2[12]) );
  degree_computation_2 degree1 ( .deg_Ri(deg_Ri), .deg_Qi(deg_Qi), .stop_i(n62), .d1out(d1out), .start(start), .deg_Ro(deg_Ro), .deg_Qo(deg_Qo), .stop_o(
        stop_o), .sw(sw), .clk(clk), .reset(reset) );
  mux_13_44 m1 ( .a(Q1), .b(R1), .sel(sw), .out(r_mux) );
  mux_13_43 m2 ( .a(R1), .b(Q1), .sel(sw), .out(q_mux) );
  mux_13_42 m3 ( .a(U1), .b(L1), .sel(sw), .out(l_mux) );
  mux_13_41 m4 ( .a(L1), .b(U1), .sel(sw), .out(u_mux) );
  feedback_ckt_11 D1 ( .Din(q_mux), .start(n2), .Qout(d1out), .clk(clk), 
        .reset(reset) );
  feedback_ckt_10 D2 ( .Din(r_mux), .start(n2), .Qout(d2out), .clk(clk), 
        .reset(reset) );
  feedback_ckt_9 D3 ( .Din(q_mux), .start(n2), .Qout(d3out), .clk(clk), 
        .reset(reset) );
  feedback_ckt_8 D4 ( .Din(r_mux), .start(n61), .Qout(d4out), .clk(clk), 
        .reset(reset) );
  multiplier_11 mx1 ( .a(R2), .b(d1out), .c(m1out) );
  multiplier_10 mx2 ( .a(d2out), .b(Q2), .c(m2out) );
  multiplier_9 mx3 ( .a(L2), .b(d3out), .c(m3out) );
  multiplier_8 mx4 ( .a(d4out), .b(U2), .c(m4out) );
  mux_13_40 m5 ( .a(R2), .b(add1out), .sel(n62), .out(Rout) );
  mux_13_39 m6 ( .a(Q2), .b(Q3), .sel(stop_i), .out(Qout) );
  mux_13_38 m7 ( .a(L2), .b(add2out), .sel(n62), .out(Lout) );
  mux_13_37 m8 ( .a(U2), .b(U3), .sel(n62), .out(Uout) );
  DFFRHQXL \R1_reg[12]  ( .D(n288), .CK(clk), .RN(reset), .Q(R1[12]) );
  DFFRHQXL \L1_reg[12]  ( .D(n345), .CK(clk), .RN(reset), .Q(L1[12]) );
  DFFRHQXL \L1_reg[2]  ( .D(n347), .CK(clk), .RN(reset), .Q(L1[2]) );
  DFFSX1 S3_reg ( .D(n402), .CK(clk), .SN(reset), .Q(st_out), .QN(n403) );
  DFFSX1 S2_reg ( .D(n287), .CK(clk), .SN(reset), .Q(S2) );
  DFFRHQX1 \Q3_reg[12]  ( .D(n332), .CK(clk), .RN(reset), .Q(Q3[12]) );
  DFFRHQX1 \Q3_reg[11]  ( .D(n333), .CK(clk), .RN(reset), .Q(Q3[11]) );
  DFFRHQX1 \Q3_reg[10]  ( .D(n334), .CK(clk), .RN(reset), .Q(Q3[10]) );
  DFFRHQX1 \Q3_reg[9]  ( .D(n335), .CK(clk), .RN(reset), .Q(Q3[9]) );
  DFFRHQX1 \Q3_reg[8]  ( .D(n336), .CK(clk), .RN(reset), .Q(Q3[8]) );
  DFFRHQX1 \Q3_reg[7]  ( .D(n337), .CK(clk), .RN(reset), .Q(Q3[7]) );
  DFFRHQX1 \Q3_reg[6]  ( .D(n338), .CK(clk), .RN(reset), .Q(Q3[6]) );
  DFFRHQX1 \Q3_reg[5]  ( .D(n339), .CK(clk), .RN(reset), .Q(Q3[5]) );
  DFFRHQX1 \Q3_reg[4]  ( .D(n340), .CK(clk), .RN(reset), .Q(Q3[4]) );
  DFFRHQX1 \Q3_reg[3]  ( .D(n341), .CK(clk), .RN(reset), .Q(Q3[3]) );
  DFFRHQX1 \Q3_reg[2]  ( .D(n342), .CK(clk), .RN(reset), .Q(Q3[2]) );
  DFFRHQX1 \Q3_reg[1]  ( .D(n343), .CK(clk), .RN(reset), .Q(Q3[1]) );
  DFFRHQX1 \Q3_reg[0]  ( .D(n344), .CK(clk), .RN(reset), .Q(Q3[0]) );
  DFFRHQX1 \U3_reg[12]  ( .D(n389), .CK(clk), .RN(reset), .Q(U3[12]) );
  DFFRHQX1 \U3_reg[11]  ( .D(n390), .CK(clk), .RN(reset), .Q(U3[11]) );
  DFFRHQX1 \U3_reg[10]  ( .D(n391), .CK(clk), .RN(reset), .Q(U3[10]) );
  DFFRHQX1 \U3_reg[9]  ( .D(n392), .CK(clk), .RN(reset), .Q(U3[9]) );
  DFFRHQX1 \U3_reg[8]  ( .D(n393), .CK(clk), .RN(reset), .Q(U3[8]) );
  DFFRHQX1 \U3_reg[7]  ( .D(n394), .CK(clk), .RN(reset), .Q(U3[7]) );
  DFFRHQX1 \U3_reg[6]  ( .D(n395), .CK(clk), .RN(reset), .Q(U3[6]) );
  DFFRHQX1 \U3_reg[5]  ( .D(n396), .CK(clk), .RN(reset), .Q(U3[5]) );
  DFFRHQX1 \U3_reg[4]  ( .D(n397), .CK(clk), .RN(reset), .Q(U3[4]) );
  DFFRHQX1 \U3_reg[3]  ( .D(n398), .CK(clk), .RN(reset), .Q(U3[3]) );
  DFFRHQX1 \U3_reg[2]  ( .D(n399), .CK(clk), .RN(reset), .Q(U3[2]) );
  DFFRHQX1 \U3_reg[1]  ( .D(n400), .CK(clk), .RN(reset), .Q(U3[1]) );
  DFFRHQX1 \U3_reg[0]  ( .D(n401), .CK(clk), .RN(reset), .Q(U3[0]) );
  DFFRHQX1 \R1_reg[6]  ( .D(n289), .CK(clk), .RN(reset), .Q(R1[6]) );
  DFFRHQX1 \R1_reg[1]  ( .D(n291), .CK(clk), .RN(reset), .Q(R1[1]) );
  DFFRHQX1 \R1_reg[0]  ( .D(n292), .CK(clk), .RN(reset), .Q(R1[0]) );
  DFFRHQX1 \Q1_reg[12]  ( .D(n293), .CK(clk), .RN(reset), .Q(Q1[12]) );
  DFFRHQX1 \Q1_reg[11]  ( .D(n294), .CK(clk), .RN(reset), .Q(Q1[11]) );
  DFFRHQX1 \Q1_reg[10]  ( .D(n295), .CK(clk), .RN(reset), .Q(Q1[10]) );
  DFFRHQX1 \Q1_reg[8]  ( .D(n297), .CK(clk), .RN(reset), .Q(Q1[8]) );
  DFFRHQX1 \Q1_reg[7]  ( .D(n298), .CK(clk), .RN(reset), .Q(Q1[7]) );
  DFFRHQX1 \Q1_reg[6]  ( .D(n299), .CK(clk), .RN(reset), .Q(Q1[6]) );
  DFFRHQX1 \Q1_reg[5]  ( .D(n300), .CK(clk), .RN(reset), .Q(Q1[5]) );
  DFFRHQX1 \Q1_reg[4]  ( .D(n301), .CK(clk), .RN(reset), .Q(Q1[4]) );
  DFFRHQX1 \Q1_reg[3]  ( .D(n302), .CK(clk), .RN(reset), .Q(Q1[3]) );
  DFFRHQX1 \Q1_reg[2]  ( .D(n303), .CK(clk), .RN(reset), .Q(Q1[2]) );
  DFFRHQX1 \Q1_reg[1]  ( .D(n304), .CK(clk), .RN(reset), .Q(Q1[1]) );
  DFFRHQX1 \Q1_reg[0]  ( .D(n305), .CK(clk), .RN(reset), .Q(Q1[0]) );
  DFFRHQX1 \L1_reg[1]  ( .D(n348), .CK(clk), .RN(reset), .Q(L1[1]) );
  DFFRHQX1 \L1_reg[0]  ( .D(n349), .CK(clk), .RN(reset), .Q(L1[0]) );
  DFFRHQX1 \U1_reg[12]  ( .D(n350), .CK(clk), .RN(reset), .Q(U1[12]) );
  DFFRHQX1 \U1_reg[11]  ( .D(n351), .CK(clk), .RN(reset), .Q(U1[11]) );
  DFFRHQX1 \U1_reg[10]  ( .D(n352), .CK(clk), .RN(reset), .Q(U1[10]) );
  DFFRHQX1 \U1_reg[8]  ( .D(n354), .CK(clk), .RN(reset), .Q(U1[8]) );
  DFFRHQX1 \U1_reg[7]  ( .D(n355), .CK(clk), .RN(reset), .Q(U1[7]) );
  DFFRHQX1 \U1_reg[6]  ( .D(n356), .CK(clk), .RN(reset), .Q(U1[6]) );
  DFFRHQX1 \U1_reg[5]  ( .D(n357), .CK(clk), .RN(reset), .Q(U1[5]) );
  DFFRHQX1 \U1_reg[4]  ( .D(n358), .CK(clk), .RN(reset), .Q(U1[4]) );
  DFFRHQX1 \U1_reg[3]  ( .D(n359), .CK(clk), .RN(reset), .Q(U1[3]) );
  DFFRHQX1 \U1_reg[2]  ( .D(n360), .CK(clk), .RN(reset), .Q(U1[2]) );
  DFFRHQX1 \U1_reg[1]  ( .D(n361), .CK(clk), .RN(reset), .Q(U1[1]) );
  DFFRHQX1 \U1_reg[0]  ( .D(n362), .CK(clk), .RN(reset), .Q(U1[0]) );
  DFFRHQX1 \Q1_reg[9]  ( .D(n296), .CK(clk), .RN(reset), .Q(Q1[9]) );
  DFFRHQX1 \U1_reg[9]  ( .D(n353), .CK(clk), .RN(reset), .Q(U1[9]) );
  DFFRHQX1 \R1_reg[11]  ( .D(n270), .CK(clk), .RN(reset), .Q(R1[11]) );
  DFFRHQX1 \R1_reg[10]  ( .D(n271), .CK(clk), .RN(reset), .Q(R1[10]) );
  DFFRHQX1 \R1_reg[8]  ( .D(n273), .CK(clk), .RN(reset), .Q(R1[8]) );
  DFFRHQX1 \R1_reg[7]  ( .D(n274), .CK(clk), .RN(reset), .Q(R1[7]) );
  DFFRHQX1 \R1_reg[5]  ( .D(n275), .CK(clk), .RN(reset), .Q(R1[5]) );
  DFFRHQX1 \R1_reg[4]  ( .D(n276), .CK(clk), .RN(reset), .Q(R1[4]) );
  DFFRHQX1 \R1_reg[3]  ( .D(n277), .CK(clk), .RN(reset), .Q(R1[3]) );
  DFFRHQX1 \L1_reg[11]  ( .D(n278), .CK(clk), .RN(reset), .Q(L1[11]) );
  DFFRHQX1 \L1_reg[10]  ( .D(n279), .CK(clk), .RN(reset), .Q(L1[10]) );
  DFFRHQX1 \L1_reg[8]  ( .D(n281), .CK(clk), .RN(reset), .Q(L1[8]) );
  DFFRHQX1 \L1_reg[7]  ( .D(n282), .CK(clk), .RN(reset), .Q(L1[7]) );
  DFFRHQX1 \L1_reg[5]  ( .D(n283), .CK(clk), .RN(reset), .Q(L1[5]) );
  DFFRHQX1 \L1_reg[4]  ( .D(n284), .CK(clk), .RN(reset), .Q(L1[4]) );
  DFFRHQX1 \L1_reg[3]  ( .D(n285), .CK(clk), .RN(reset), .Q(L1[3]) );
  DFFRHQX1 \R1_reg[9]  ( .D(n272), .CK(clk), .RN(reset), .Q(R1[9]) );
  DFFRHQX1 \L1_reg[9]  ( .D(n280), .CK(clk), .RN(reset), .Q(L1[9]) );
  DFFSX1 S1_reg ( .D(n286), .CK(clk), .SN(reset), .Q(n2), .QN(n57) );
  DFFRHQX1 \L2_reg[0]  ( .D(n376), .CK(clk), .RN(reset), .Q(L2[0]) );
  DFFRHQX1 \R2_reg[0]  ( .D(n319), .CK(clk), .RN(reset), .Q(R2[0]) );
  DFFRHQX1 \R2_reg[1]  ( .D(n320), .CK(clk), .RN(reset), .Q(R2[1]) );
  DFFRHQX1 \R2_reg[2]  ( .D(n321), .CK(clk), .RN(reset), .Q(R2[2]) );
  DFFRHQX1 \R2_reg[6]  ( .D(n325), .CK(clk), .RN(reset), .Q(R2[6]) );
  DFFRHQX1 \L2_reg[1]  ( .D(n377), .CK(clk), .RN(reset), .Q(L2[1]) );
  DFFRHQX1 \L2_reg[2]  ( .D(n378), .CK(clk), .RN(reset), .Q(L2[2]) );
  DFFRHQX1 \L2_reg[6]  ( .D(n382), .CK(clk), .RN(reset), .Q(L2[6]) );
  DFFRHQX1 \R2_reg[3]  ( .D(n322), .CK(clk), .RN(reset), .Q(R2[3]) );
  DFFRHQX1 \R2_reg[4]  ( .D(n323), .CK(clk), .RN(reset), .Q(R2[4]) );
  DFFRHQX1 \R2_reg[5]  ( .D(n324), .CK(clk), .RN(reset), .Q(R2[5]) );
  DFFRHQX1 \R2_reg[7]  ( .D(n326), .CK(clk), .RN(reset), .Q(R2[7]) );
  DFFRHQX1 \R2_reg[8]  ( .D(n327), .CK(clk), .RN(reset), .Q(R2[8]) );
  DFFRHQX1 \R2_reg[9]  ( .D(n328), .CK(clk), .RN(reset), .Q(R2[9]) );
  DFFRHQX1 \R2_reg[10]  ( .D(n329), .CK(clk), .RN(reset), .Q(R2[10]) );
  DFFRHQX1 \L2_reg[3]  ( .D(n379), .CK(clk), .RN(reset), .Q(L2[3]) );
  DFFRHQX1 \L2_reg[4]  ( .D(n380), .CK(clk), .RN(reset), .Q(L2[4]) );
  DFFRHQX1 \L2_reg[5]  ( .D(n381), .CK(clk), .RN(reset), .Q(L2[5]) );
  DFFRHQX1 \L2_reg[7]  ( .D(n383), .CK(clk), .RN(reset), .Q(L2[7]) );
  DFFRHQX1 \L2_reg[8]  ( .D(n384), .CK(clk), .RN(reset), .Q(L2[8]) );
  DFFRHQX1 \L2_reg[9]  ( .D(n385), .CK(clk), .RN(reset), .Q(L2[9]) );
  DFFRHQX1 \L2_reg[10]  ( .D(n386), .CK(clk), .RN(reset), .Q(L2[10]) );
  DFFRHQX1 \Q2_reg[2]  ( .D(n308), .CK(clk), .RN(reset), .Q(Q2[2]) );
  DFFRHQX1 \Q2_reg[5]  ( .D(n311), .CK(clk), .RN(reset), .Q(Q2[5]) );
  DFFRHQX1 \Q2_reg[6]  ( .D(n312), .CK(clk), .RN(reset), .Q(Q2[6]) );
  DFFRHQX1 \Q2_reg[7]  ( .D(n313), .CK(clk), .RN(reset), .Q(Q2[7]) );
  DFFRHQX1 \Q2_reg[8]  ( .D(n314), .CK(clk), .RN(reset), .Q(Q2[8]) );
  DFFRHQX1 \Q2_reg[12]  ( .D(n318), .CK(clk), .RN(reset), .Q(Q2[12]) );
  DFFRHQX1 \U2_reg[2]  ( .D(n365), .CK(clk), .RN(reset), .Q(U2[2]) );
  DFFRHQX1 \U2_reg[5]  ( .D(n368), .CK(clk), .RN(reset), .Q(U2[5]) );
  DFFRHQX1 \U2_reg[6]  ( .D(n369), .CK(clk), .RN(reset), .Q(U2[6]) );
  DFFRHQX1 \U2_reg[7]  ( .D(n370), .CK(clk), .RN(reset), .Q(U2[7]) );
  DFFRHQX1 \U2_reg[8]  ( .D(n371), .CK(clk), .RN(reset), .Q(U2[8]) );
  DFFRHQX1 \U2_reg[12]  ( .D(n375), .CK(clk), .RN(reset), .Q(U2[12]) );
  DFFRHQX1 \Q2_reg[9]  ( .D(n315), .CK(clk), .RN(reset), .Q(Q2[9]) );
  DFFRHQX1 \U2_reg[9]  ( .D(n372), .CK(clk), .RN(reset), .Q(U2[9]) );
  DFFRHQX1 \Q2_reg[0]  ( .D(n306), .CK(clk), .RN(reset), .Q(Q2[0]) );
  DFFRHQX1 \U2_reg[0]  ( .D(n363), .CK(clk), .RN(reset), .Q(U2[0]) );
  DFFRHQX1 \Q2_reg[1]  ( .D(n307), .CK(clk), .RN(reset), .Q(Q2[1]) );
  DFFRHQX1 \U2_reg[1]  ( .D(n364), .CK(clk), .RN(reset), .Q(U2[1]) );
  DFFRHQX2 \U2_reg[11]  ( .D(n374), .CK(clk), .RN(reset), .Q(U2[11]) );
  DFFRHQX2 \Q2_reg[4]  ( .D(n310), .CK(clk), .RN(reset), .Q(Q2[4]) );
  DFFRHQX2 \U2_reg[4]  ( .D(n367), .CK(clk), .RN(reset), .Q(U2[4]) );
  DFFRHQX2 \U2_reg[10]  ( .D(n373), .CK(clk), .RN(reset), .Q(U2[10]) );
  DFFRHQX2 \L2_reg[11]  ( .D(n387), .CK(clk), .RN(reset), .Q(L2[11]) );
  DFFRHQXL \R1_reg[2]  ( .D(n290), .CK(clk), .RN(reset), .Q(R1[2]) );
  DFFRHQX2 \Q2_reg[3]  ( .D(n309), .CK(clk), .RN(reset), .Q(Q2[3]) );
  DFFRHQX2 \Q2_reg[10]  ( .D(n316), .CK(clk), .RN(reset), .Q(Q2[10]) );
  DFFRHQX2 \U2_reg[3]  ( .D(n366), .CK(clk), .RN(reset), .Q(U2[3]) );
  DFFRHQXL \L1_reg[6]  ( .D(n346), .CK(clk), .RN(reset), .Q(L1[6]) );
  DFFRHQX2 \Q2_reg[11]  ( .D(n317), .CK(clk), .RN(reset), .Q(Q2[11]) );
  DFFRHQX2 \R2_reg[11]  ( .D(n330), .CK(clk), .RN(reset), .Q(R2[11]) );
  MX2X2 U2_inst ( .A(R1[5]), .B(Rin[5]), .S0(n264), .Y(n275) );
  MX2X1 U3_inst ( .A(R1[8]), .B(Rin[8]), .S0(n201), .Y(n273) );
  INVX1 U4 ( .A(L1[12]), .Y(n58) );
  AOI22XL U5 ( .A0(n122), .A1(U2[2]), .B0(U3[2]), .B1(n65), .Y(n517) );
  AOI22X1 U6 ( .A0(Rin[12]), .A1(n64), .B0(R1[12]), .B1(n134), .Y(n406) );
  MX2X2 U7 ( .A(L1[5]), .B(Lin[5]), .S0(n200), .Y(n283) );
  AOI2BB2X1 U8 ( .B0(Lin[12]), .B1(n263), .A0N(n58), .A1N(n258), .Y(n463) );
  MX2X1 U9 ( .A(L1[8]), .B(Lin[8]), .S0(n195), .Y(n281) );
  MX2X1 U10 ( .A(R1[3]), .B(Rin[3]), .S0(n262), .Y(n277) );
  MX2X1 U11 ( .A(R1[10]), .B(Rin[10]), .S0(n265), .Y(n271) );
  MX2X1 U12 ( .A(L1[10]), .B(Lin[10]), .S0(start_cnt), .Y(n279) );
  MX2X1 U13 ( .A(L1[3]), .B(Lin[3]), .S0(n259), .Y(n285) );
  MX2X1 U14 ( .A(L1[11]), .B(Lin[11]), .S0(n265), .Y(n278) );
  MX2X1 U15 ( .A(R1[4]), .B(Rin[4]), .S0(n197), .Y(n276) );
  MX2X1 U16 ( .A(L1[7]), .B(Lin[7]), .S0(n198), .Y(n282) );
  MX2X1 U17 ( .A(L1[4]), .B(Lin[4]), .S0(n195), .Y(n284) );
  MX2X1 U18 ( .A(R1[11]), .B(Rin[11]), .S0(n265), .Y(n270) );
  MX2X1 U19 ( .A(R1[7]), .B(Rin[7]), .S0(n260), .Y(n274) );
  XOR2X1 U20 ( .A(m2out[4]), .B(m1out[4]), .Y(add1out[4]) );
  XOR2X1 U21 ( .A(m4out[8]), .B(m3out[8]), .Y(add2out[8]) );
  XOR2X1 U22 ( .A(m4out[11]), .B(m3out[11]), .Y(add2out[11]) );
  XOR2X1 U23 ( .A(m4out[5]), .B(m3out[5]), .Y(add2out[5]) );
  XOR2X1 U24 ( .A(m2out[5]), .B(m1out[5]), .Y(add1out[5]) );
  MX2X1 U25 ( .A(L1[9]), .B(Lin[9]), .S0(n64), .Y(n280) );
  MX2X1 U26 ( .A(R1[9]), .B(Rin[9]), .S0(n258), .Y(n272) );
  INVXL U27 ( .A(n406), .Y(n288) );
  INVXL U28 ( .A(n463), .Y(n345) );
  INVXL U29 ( .A(n465), .Y(n347) );
  INVXL U30 ( .A(n407), .Y(n289) );
  INVXL U31 ( .A(n409), .Y(n291) );
  INVXL U32 ( .A(n408), .Y(n290) );
  INVXL U33 ( .A(n464), .Y(n346) );
  INVXL U34 ( .A(n466), .Y(n348) );
  AOI22XL U35 ( .A0(n262), .A1(Q2[1]), .B0(Q3[1]), .B1(n123), .Y(n461) );
  AOI22XL U36 ( .A0(L2[12]), .A1(n193), .B0(l_mux[12]), .B1(n264), .Y(n506) );
  AOI22XL U37 ( .A0(n194), .A1(U2[11]), .B0(u_mux[11]), .B1(n263), .Y(n492) );
  AOI22XL U38 ( .A0(n128), .A1(U2[10]), .B0(u_mux[10]), .B1(n197), .Y(n491) );
  AOI22XL U39 ( .A0(n134), .A1(U2[3]), .B0(u_mux[3]), .B1(n265), .Y(n484) );
  AOI22XL U40 ( .A0(R2[12]), .A1(n128), .B0(r_mux[12]), .B1(n259), .Y(n449) );
  AOI22XL U41 ( .A0(R2[11]), .A1(n124), .B0(r_mux[11]), .B1(n262), .Y(n448) );
  AOI22XL U42 ( .A0(n124), .A1(Q2[11]), .B0(q_mux[11]), .B1(n260), .Y(n435) );
  AOI22XL U43 ( .A0(n124), .A1(Q2[3]), .B0(q_mux[3]), .B1(n198), .Y(n427) );
  AOI22XL U44 ( .A0(n262), .A1(U2[0]), .B0(U3[0]), .B1(n65), .Y(n519) );
  AOI22XL U45 ( .A0(n200), .A1(U2[1]), .B0(U3[1]), .B1(n266), .Y(n518) );
  AOI22XL U46 ( .A0(L2[9]), .A1(n193), .B0(l_mux[9]), .B1(n265), .Y(n503) );
  AOI22XL U47 ( .A0(L2[8]), .A1(n136), .B0(l_mux[8]), .B1(n259), .Y(n502) );
  AOI22XL U48 ( .A0(L2[5]), .A1(n136), .B0(l_mux[5]), .B1(n199), .Y(n499) );
  AOI22XL U49 ( .A0(L2[3]), .A1(n128), .B0(l_mux[3]), .B1(n201), .Y(n497) );
  AOI22XL U50 ( .A0(n130), .A1(U2[12]), .B0(u_mux[12]), .B1(n263), .Y(n493) );
  AOI22XL U51 ( .A0(n193), .A1(U2[9]), .B0(u_mux[9]), .B1(n262), .Y(n490) );
  AOI22XL U52 ( .A0(n129), .A1(U2[8]), .B0(u_mux[8]), .B1(n258), .Y(n489) );
  AOI22XL U53 ( .A0(n193), .A1(U2[7]), .B0(u_mux[7]), .B1(n195), .Y(n488) );
  AOI22XL U54 ( .A0(n136), .A1(U2[6]), .B0(u_mux[6]), .B1(n197), .Y(n487) );
  AOI22XL U55 ( .A0(n136), .A1(U2[5]), .B0(u_mux[5]), .B1(n258), .Y(n486) );
  AOI22XL U56 ( .A0(n127), .A1(U2[4]), .B0(u_mux[4]), .B1(n195), .Y(n485) );
  AOI22XL U57 ( .A0(n130), .A1(U2[1]), .B0(u_mux[1]), .B1(n199), .Y(n482) );
  AOI22XL U58 ( .A0(n128), .A1(U2[0]), .B0(u_mux[0]), .B1(n264), .Y(n481) );
  AOI22XL U59 ( .A0(R2[10]), .A1(n128), .B0(r_mux[10]), .B1(n258), .Y(n447) );
  AOI22XL U60 ( .A0(R2[9]), .A1(n124), .B0(r_mux[9]), .B1(n200), .Y(n446) );
  AOI22XL U61 ( .A0(R2[8]), .A1(n128), .B0(r_mux[8]), .B1(n201), .Y(n445) );
  AOI22XL U62 ( .A0(R2[7]), .A1(n134), .B0(r_mux[7]), .B1(n262), .Y(n444) );
  AOI22XL U63 ( .A0(R2[6]), .A1(n130), .B0(r_mux[6]), .B1(n198), .Y(n443) );
  AOI22XL U64 ( .A0(R2[5]), .A1(n126), .B0(r_mux[5]), .B1(n260), .Y(n442) );
  AOI22XL U65 ( .A0(R2[4]), .A1(n130), .B0(r_mux[4]), .B1(n259), .Y(n441) );
  AOI22XL U66 ( .A0(R2[3]), .A1(n65), .B0(r_mux[3]), .B1(n259), .Y(n440) );
  AOI22XL U67 ( .A0(n128), .A1(Q2[12]), .B0(q_mux[12]), .B1(n195), .Y(n436) );
  AOI22XL U68 ( .A0(n123), .A1(Q2[9]), .B0(q_mux[9]), .B1(n200), .Y(n433) );
  AOI22XL U69 ( .A0(n126), .A1(Q2[8]), .B0(q_mux[8]), .B1(n64), .Y(n432) );
  AOI22XL U70 ( .A0(n124), .A1(Q2[7]), .B0(q_mux[7]), .B1(n262), .Y(n431) );
  AOI22XL U71 ( .A0(n128), .A1(Q2[6]), .B0(q_mux[6]), .B1(n201), .Y(n430) );
  AOI22XL U72 ( .A0(n123), .A1(Q2[5]), .B0(q_mux[5]), .B1(n197), .Y(n429) );
  AOI22XL U73 ( .A0(n194), .A1(Q2[4]), .B0(q_mux[4]), .B1(n199), .Y(n428) );
  AOI22XL U74 ( .A0(n126), .A1(Q2[2]), .B0(q_mux[2]), .B1(n199), .Y(n426) );
  AOI22XL U75 ( .A0(n123), .A1(Q2[1]), .B0(q_mux[1]), .B1(n265), .Y(n425) );
  AOI22XL U76 ( .A0(n123), .A1(Q2[0]), .B0(q_mux[0]), .B1(n64), .Y(n424) );
  AOI22XL U77 ( .A0(n122), .A1(U2[3]), .B0(U3[3]), .B1(n65), .Y(n516) );
  AOI22XL U78 ( .A0(n122), .A1(U2[4]), .B0(U3[4]), .B1(n266), .Y(n515) );
  AOI22XL U79 ( .A0(n122), .A1(U2[5]), .B0(U3[5]), .B1(n126), .Y(n514) );
  AOI22XL U80 ( .A0(n122), .A1(U2[6]), .B0(U3[6]), .B1(n127), .Y(n513) );
  AOI22XL U81 ( .A0(n122), .A1(U2[7]), .B0(U3[7]), .B1(n193), .Y(n512) );
  AOI22XL U82 ( .A0(n122), .A1(U2[8]), .B0(U3[8]), .B1(n136), .Y(n511) );
  AOI22XL U83 ( .A0(n122), .A1(U2[9]), .B0(U3[9]), .B1(n129), .Y(n510) );
  AOI22XL U84 ( .A0(n122), .A1(U2[10]), .B0(U3[10]), .B1(n134), .Y(n509) );
  AOI22XL U85 ( .A0(n122), .A1(U2[11]), .B0(U3[11]), .B1(n126), .Y(n508) );
  AOI22XL U86 ( .A0(n265), .A1(U2[12]), .B0(U3[12]), .B1(n130), .Y(n507) );
  AOI22XL U87 ( .A0(n64), .A1(Q2[0]), .B0(Q3[0]), .B1(n127), .Y(n462) );
  AOI22XL U88 ( .A0(n197), .A1(Q2[2]), .B0(Q3[2]), .B1(n65), .Y(n460) );
  AOI22XL U89 ( .A0(n198), .A1(Q2[3]), .B0(Q3[3]), .B1(n194), .Y(n459) );
  AOI22XL U90 ( .A0(n263), .A1(Q2[4]), .B0(Q3[4]), .B1(n266), .Y(n458) );
  AOI22XL U91 ( .A0(n64), .A1(Q2[5]), .B0(Q3[5]), .B1(n194), .Y(n457) );
  AOI22XL U92 ( .A0(n260), .A1(Q2[6]), .B0(Q3[6]), .B1(n127), .Y(n456) );
  AOI22XL U93 ( .A0(n264), .A1(Q2[9]), .B0(Q3[9]), .B1(n266), .Y(n453) );
  AOI22XL U94 ( .A0(n195), .A1(Q2[12]), .B0(Q3[12]), .B1(n130), .Y(n450) );
  AOI22XL U95 ( .A0(n195), .A1(Q2[7]), .B0(Q3[7]), .B1(n130), .Y(n455) );
  AOI22XL U96 ( .A0(n200), .A1(Q2[8]), .B0(Q3[8]), .B1(n266), .Y(n454) );
  AOI22XL U97 ( .A0(n259), .A1(Q2[11]), .B0(Q3[11]), .B1(n65), .Y(n451) );
  AOI22XL U98 ( .A0(L2[11]), .A1(n134), .B0(l_mux[11]), .B1(n201), .Y(n505) );
  AOI22XL U99 ( .A0(L2[10]), .A1(n127), .B0(l_mux[10]), .B1(n265), .Y(n504) );
  INVX1 U100 ( .A(n129), .Y(n122) );
  INVX1 U101 ( .A(n201), .Y(n123) );
  INVX1 U102 ( .A(n200), .Y(n124) );
  INVX1 U103 ( .A(n197), .Y(n193) );
  INVX1 U104 ( .A(n197), .Y(n136) );
  INVX1 U105 ( .A(n198), .Y(n134) );
  INVX1 U106 ( .A(n198), .Y(n130) );
  INVX1 U107 ( .A(n199), .Y(n128) );
  INVX1 U108 ( .A(n199), .Y(n127) );
  INVX1 U109 ( .A(n199), .Y(n126) );
  INVX1 U110 ( .A(n198), .Y(n129) );
  INVX1 U111 ( .A(n197), .Y(n194) );
  INVX1 U112 ( .A(n127), .Y(n201) );
  INVX1 U113 ( .A(n266), .Y(n197) );
  INVX1 U114 ( .A(n266), .Y(n195) );
  INVX1 U115 ( .A(n136), .Y(n258) );
  INVX1 U116 ( .A(n134), .Y(n262) );
  INVX1 U117 ( .A(n65), .Y(n259) );
  INVX1 U118 ( .A(n193), .Y(n260) );
  INVX1 U119 ( .A(n266), .Y(n199) );
  INVX1 U120 ( .A(n194), .Y(n200) );
  INVX1 U121 ( .A(n266), .Y(n263) );
  INVX1 U122 ( .A(n65), .Y(n264) );
  INVX1 U123 ( .A(n65), .Y(n265) );
  INVX1 U124 ( .A(n266), .Y(n198) );
  INVX1 U125 ( .A(n64), .Y(n266) );
  INVX1 U126 ( .A(n65), .Y(n64) );
  INVX1 U127 ( .A(start_cnt), .Y(n65) );
  XOR2X1 U128 ( .A(m3out[10]), .B(m4out[10]), .Y(add2out[10]) );
  XOR2X1 U129 ( .A(m1out[10]), .B(m2out[10]), .Y(add1out[10]) );
  XOR2X1 U130 ( .A(m1out[8]), .B(m2out[8]), .Y(add1out[8]) );
  XOR2X1 U131 ( .A(m4out[6]), .B(m3out[6]), .Y(add2out[6]) );
  XOR2X1 U132 ( .A(m2out[6]), .B(m1out[6]), .Y(add1out[6]) );
  XOR2X1 U133 ( .A(m2out[2]), .B(m1out[2]), .Y(add1out[2]) );
  XOR2X1 U134 ( .A(m4out[1]), .B(m3out[1]), .Y(add2out[1]) );
  XOR2X1 U135 ( .A(m4out[2]), .B(m3out[2]), .Y(add2out[2]) );
  XOR2X1 U136 ( .A(m2out[1]), .B(m1out[1]), .Y(add1out[1]) );
  XOR2X1 U137 ( .A(m4out[12]), .B(m3out[12]), .Y(add2out[12]) );
  XOR2X1 U138 ( .A(m2out[12]), .B(m1out[12]), .Y(add1out[12]) );
  XOR2X1 U139 ( .A(m1out[7]), .B(m2out[7]), .Y(add1out[7]) );
  XOR2X1 U140 ( .A(m3out[7]), .B(m4out[7]), .Y(add2out[7]) );
  XOR2X1 U141 ( .A(m3out[3]), .B(m4out[3]), .Y(add2out[3]) );
  XOR2X1 U142 ( .A(m3out[4]), .B(m4out[4]), .Y(add2out[4]) );
  XOR2X1 U143 ( .A(m3out[9]), .B(m4out[9]), .Y(add2out[9]) );
  XOR2X1 U144 ( .A(m1out[3]), .B(m2out[3]), .Y(add1out[3]) );
  XOR2X1 U145 ( .A(m1out[9]), .B(m2out[9]), .Y(add1out[9]) );
  XOR2X1 U146 ( .A(m1out[11]), .B(m2out[11]), .Y(add1out[11]) );
  XOR2X1 U147 ( .A(m2out[0]), .B(m1out[0]), .Y(add1out[0]) );
  XOR2X1 U148 ( .A(m4out[0]), .B(m3out[0]), .Y(add2out[0]) );
  INVX1 U149 ( .A(n57), .Y(n61) );
  INVX1 U150 ( .A(n63), .Y(n62) );
  OAI2BB2X1 U151 ( .B0(n198), .B1(n403), .A0N(S2), .A1N(n263), .Y(n402) );
  AOI22X1 U152 ( .A0(L1[2]), .A1(n126), .B0(Lin[2]), .B1(n199), .Y(n465) );
  INVX1 U153 ( .A(n518), .Y(n400) );
  INVX1 U154 ( .A(n482), .Y(n364) );
  INVX1 U155 ( .A(n461), .Y(n343) );
  INVX1 U156 ( .A(n425), .Y(n307) );
  INVX1 U157 ( .A(n519), .Y(n401) );
  INVX1 U158 ( .A(n481), .Y(n363) );
  INVX1 U159 ( .A(n462), .Y(n344) );
  INVX1 U160 ( .A(n424), .Y(n306) );
  INVX1 U161 ( .A(n510), .Y(n392) );
  INVX1 U162 ( .A(n490), .Y(n372) );
  INVX1 U163 ( .A(n453), .Y(n335) );
  INVX1 U164 ( .A(n433), .Y(n315) );
  INVX1 U165 ( .A(n517), .Y(n399) );
  INVX1 U166 ( .A(n516), .Y(n398) );
  INVX1 U167 ( .A(n515), .Y(n397) );
  INVX1 U168 ( .A(n514), .Y(n396) );
  INVX1 U169 ( .A(n513), .Y(n395) );
  INVX1 U170 ( .A(n512), .Y(n394) );
  INVX1 U171 ( .A(n511), .Y(n393) );
  INVX1 U172 ( .A(n509), .Y(n391) );
  INVX1 U173 ( .A(n508), .Y(n390) );
  INVX1 U174 ( .A(n507), .Y(n389) );
  INVX1 U175 ( .A(n493), .Y(n375) );
  INVX1 U176 ( .A(n492), .Y(n374) );
  INVX1 U177 ( .A(n491), .Y(n373) );
  INVX1 U178 ( .A(n489), .Y(n371) );
  INVX1 U179 ( .A(n488), .Y(n370) );
  INVX1 U180 ( .A(n487), .Y(n369) );
  INVX1 U181 ( .A(n486), .Y(n368) );
  INVX1 U182 ( .A(n485), .Y(n367) );
  INVX1 U183 ( .A(n484), .Y(n366) );
  INVX1 U184 ( .A(n483), .Y(n365) );
  AOI22X1 U185 ( .A0(n134), .A1(U2[2]), .B0(u_mux[2]), .B1(n200), .Y(n483) );
  INVX1 U186 ( .A(n460), .Y(n342) );
  INVX1 U187 ( .A(n459), .Y(n341) );
  INVX1 U188 ( .A(n458), .Y(n340) );
  INVX1 U189 ( .A(n457), .Y(n339) );
  INVX1 U190 ( .A(n456), .Y(n338) );
  INVX1 U191 ( .A(n455), .Y(n337) );
  INVX1 U192 ( .A(n454), .Y(n336) );
  INVX1 U193 ( .A(n452), .Y(n334) );
  AOI22X1 U194 ( .A0(n258), .A1(Q2[10]), .B0(Q3[10]), .B1(n130), .Y(n452) );
  INVX1 U195 ( .A(n450), .Y(n332) );
  INVX1 U196 ( .A(n436), .Y(n318) );
  INVX1 U197 ( .A(n434), .Y(n316) );
  AOI22X1 U198 ( .A0(n127), .A1(Q2[10]), .B0(q_mux[10]), .B1(n260), .Y(n434)
         );
  INVX1 U199 ( .A(n432), .Y(n314) );
  INVX1 U200 ( .A(n431), .Y(n313) );
  INVX1 U201 ( .A(n430), .Y(n312) );
  INVX1 U202 ( .A(n429), .Y(n311) );
  INVX1 U203 ( .A(n428), .Y(n310) );
  INVX1 U204 ( .A(n427), .Y(n309) );
  INVX1 U205 ( .A(n426), .Y(n308) );
  INVX1 U206 ( .A(n451), .Y(n333) );
  INVX1 U207 ( .A(n435), .Y(n317) );
  INVX1 U208 ( .A(n480), .Y(n362) );
  AOI22X1 U209 ( .A0(U1[0]), .A1(n124), .B0(Uin[0]), .B1(n201), .Y(n480) );
  INVX1 U210 ( .A(n479), .Y(n361) );
  AOI22X1 U211 ( .A0(U1[1]), .A1(n136), .B0(Uin[1]), .B1(n198), .Y(n479) );
  INVX1 U212 ( .A(n478), .Y(n360) );
  AOI22X1 U213 ( .A0(U1[2]), .A1(n136), .B0(Uin[2]), .B1(n199), .Y(n478) );
  INVX1 U214 ( .A(n477), .Y(n359) );
  AOI22X1 U215 ( .A0(U1[3]), .A1(n129), .B0(Uin[3]), .B1(n195), .Y(n477) );
  INVX1 U216 ( .A(n476), .Y(n358) );
  AOI22X1 U217 ( .A0(U1[4]), .A1(n126), .B0(Uin[4]), .B1(n263), .Y(n476) );
  INVX1 U218 ( .A(n475), .Y(n357) );
  AOI22X1 U219 ( .A0(U1[5]), .A1(n128), .B0(Uin[5]), .B1(n258), .Y(n475) );
  INVX1 U220 ( .A(n474), .Y(n356) );
  AOI22X1 U221 ( .A0(U1[6]), .A1(n124), .B0(Uin[6]), .B1(start_cnt), .Y(n474)
         );
  INVX1 U222 ( .A(n503), .Y(n385) );
  INVX1 U223 ( .A(n502), .Y(n384) );
  INVX1 U224 ( .A(n501), .Y(n383) );
  AOI22X1 U225 ( .A0(L2[7]), .A1(n193), .B0(l_mux[7]), .B1(n64), .Y(n501) );
  INVX1 U226 ( .A(n500), .Y(n382) );
  AOI22X1 U227 ( .A0(L2[6]), .A1(n194), .B0(l_mux[6]), .B1(n197), .Y(n500) );
  INVX1 U228 ( .A(n499), .Y(n381) );
  INVX1 U229 ( .A(n498), .Y(n380) );
  AOI22X1 U230 ( .A0(L2[4]), .A1(n130), .B0(l_mux[4]), .B1(n195), .Y(n498) );
  INVX1 U231 ( .A(n497), .Y(n379) );
  INVX1 U232 ( .A(n496), .Y(n378) );
  AOI22X1 U233 ( .A0(L2[2]), .A1(n127), .B0(l_mux[2]), .B1(n263), .Y(n496) );
  INVX1 U234 ( .A(n495), .Y(n377) );
  AOI22X1 U235 ( .A0(L2[1]), .A1(n126), .B0(l_mux[1]), .B1(n201), .Y(n495) );
  INVX1 U236 ( .A(n494), .Y(n376) );
  AOI22X1 U237 ( .A0(L2[0]), .A1(n129), .B0(l_mux[0]), .B1(n264), .Y(n494) );
  INVX1 U238 ( .A(n473), .Y(n355) );
  AOI22X1 U239 ( .A0(U1[7]), .A1(n136), .B0(Uin[7]), .B1(n260), .Y(n473) );
  INVX1 U240 ( .A(n472), .Y(n354) );
  AOI22X1 U241 ( .A0(U1[8]), .A1(n123), .B0(Uin[8]), .B1(n262), .Y(n472) );
  INVX1 U242 ( .A(n471), .Y(n353) );
  AOI22X1 U243 ( .A0(U1[9]), .A1(n130), .B0(Uin[9]), .B1(n264), .Y(n471) );
  INVX1 U244 ( .A(n470), .Y(n352) );
  AOI22X1 U245 ( .A0(U1[10]), .A1(n124), .B0(Uin[10]), .B1(n258), .Y(n470) );
  INVX1 U246 ( .A(n469), .Y(n351) );
  AOI22X1 U247 ( .A0(U1[11]), .A1(n127), .B0(Uin[11]), .B1(n195), .Y(n469) );
  INVX1 U248 ( .A(n468), .Y(n350) );
  AOI22X1 U249 ( .A0(U1[12]), .A1(n127), .B0(Uin[12]), .B1(n197), .Y(n468) );
  INVX1 U250 ( .A(n467), .Y(n349) );
  AOI22X1 U251 ( .A0(L1[0]), .A1(n128), .B0(Lin[0]), .B1(n259), .Y(n467) );
  AOI22X1 U252 ( .A0(L1[1]), .A1(n123), .B0(Lin[1]), .B1(n260), .Y(n466) );
  AOI22X1 U253 ( .A0(L1[6]), .A1(n123), .B0(Lin[6]), .B1(n200), .Y(n464) );
  INVX1 U254 ( .A(n449), .Y(n331) );
  INVX1 U255 ( .A(n448), .Y(n330) );
  INVX1 U256 ( .A(n447), .Y(n329) );
  INVX1 U257 ( .A(n446), .Y(n328) );
  INVX1 U258 ( .A(n445), .Y(n327) );
  INVX1 U259 ( .A(n444), .Y(n326) );
  INVX1 U260 ( .A(n443), .Y(n325) );
  INVX1 U261 ( .A(n442), .Y(n324) );
  INVX1 U262 ( .A(n441), .Y(n323) );
  INVX1 U263 ( .A(n440), .Y(n322) );
  INVX1 U264 ( .A(n439), .Y(n321) );
  AOI22X1 U265 ( .A0(R2[2]), .A1(n194), .B0(r_mux[2]), .B1(n198), .Y(n439) );
  INVX1 U266 ( .A(n438), .Y(n320) );
  AOI22X1 U267 ( .A0(R2[1]), .A1(n134), .B0(r_mux[1]), .B1(n265), .Y(n438) );
  INVX1 U268 ( .A(n437), .Y(n319) );
  AOI22X1 U269 ( .A0(R2[0]), .A1(n126), .B0(r_mux[0]), .B1(n263), .Y(n437) );
  INVX1 U270 ( .A(n423), .Y(n305) );
  AOI22X1 U271 ( .A0(Q1[0]), .A1(n129), .B0(Qin[0]), .B1(start_cnt), .Y(n423)
         );
  INVX1 U272 ( .A(n422), .Y(n304) );
  AOI22X1 U273 ( .A0(Q1[1]), .A1(n123), .B0(Qin[1]), .B1(n263), .Y(n422) );
  INVX1 U274 ( .A(n421), .Y(n303) );
  AOI22X1 U275 ( .A0(Q1[2]), .A1(n194), .B0(Qin[2]), .B1(n260), .Y(n421) );
  INVX1 U276 ( .A(n420), .Y(n302) );
  AOI22X1 U277 ( .A0(Q1[3]), .A1(n193), .B0(Qin[3]), .B1(start_cnt), .Y(n420)
         );
  INVX1 U278 ( .A(n419), .Y(n301) );
  AOI22X1 U279 ( .A0(Q1[4]), .A1(n194), .B0(Qin[4]), .B1(start_cnt), .Y(n419)
         );
  INVX1 U280 ( .A(n418), .Y(n300) );
  AOI22X1 U281 ( .A0(Q1[5]), .A1(n124), .B0(Qin[5]), .B1(n260), .Y(n418) );
  INVX1 U282 ( .A(n417), .Y(n299) );
  AOI22X1 U283 ( .A0(Q1[6]), .A1(n136), .B0(Qin[6]), .B1(n258), .Y(n417) );
  INVX1 U284 ( .A(n416), .Y(n298) );
  AOI22X1 U285 ( .A0(Q1[7]), .A1(n134), .B0(Qin[7]), .B1(start_cnt), .Y(n416)
         );
  INVX1 U286 ( .A(n415), .Y(n297) );
  AOI22X1 U287 ( .A0(Q1[8]), .A1(n134), .B0(Qin[8]), .B1(n258), .Y(n415) );
  INVX1 U288 ( .A(n414), .Y(n296) );
  AOI22X1 U289 ( .A0(Q1[9]), .A1(n129), .B0(Qin[9]), .B1(n265), .Y(n414) );
  INVX1 U290 ( .A(n413), .Y(n295) );
  AOI22X1 U291 ( .A0(Q1[10]), .A1(n129), .B0(Qin[10]), .B1(n262), .Y(n413) );
  INVX1 U292 ( .A(n412), .Y(n294) );
  AOI22X1 U293 ( .A0(Q1[11]), .A1(n193), .B0(Qin[11]), .B1(n259), .Y(n412) );
  INVX1 U294 ( .A(n411), .Y(n293) );
  AOI22X1 U295 ( .A0(Q1[12]), .A1(n124), .B0(Qin[12]), .B1(n262), .Y(n411) );
  INVX1 U296 ( .A(n410), .Y(n292) );
  AOI22X1 U297 ( .A0(R1[0]), .A1(n126), .B0(Rin[0]), .B1(n259), .Y(n410) );
  AOI22X1 U298 ( .A0(R1[1]), .A1(n129), .B0(Rin[1]), .B1(n264), .Y(n409) );
  AOI22X1 U299 ( .A0(R1[6]), .A1(n194), .B0(Rin[6]), .B1(n263), .Y(n407) );
  INVX1 U300 ( .A(n506), .Y(n388) );
  INVX1 U301 ( .A(n505), .Y(n387) );
  INVX1 U302 ( .A(n504), .Y(n386) );
  AOI22X1 U303 ( .A0(R1[2]), .A1(n123), .B0(Rin[2]), .B1(n260), .Y(n408) );
  INVX1 U304 ( .A(n404), .Y(n286) );
  AOI22X1 U305 ( .A0(n129), .A1(n61), .B0(start), .B1(n264), .Y(n404) );
  INVX1 U306 ( .A(n405), .Y(n287) );
  AOI22X1 U307 ( .A0(n199), .A1(n61), .B0(n193), .B1(S2), .Y(n405) );
  INVX1 U308 ( .A(stop_i), .Y(n63) );
endmodule


module euclidean_cell_1 ( deg_Ri, deg_Qi, stop_i, Rin, Qin, Lin, Uin, start, 
        start_cnt, deg_Ro, deg_Qo, stop_o, Rout, Qout, Lout, Uout, st_out, clk, 
        reset );
  input [4:0] deg_Ri;
  input [4:0] deg_Qi;
  input [12:0] Rin;
  input [12:0] Qin;
  input [12:0] Lin;
  input [12:0] Uin;
  output [4:0] deg_Ro;
  output [4:0] deg_Qo;
  output [12:0] Rout;
  output [12:0] Qout;
  output [12:0] Lout;
  output [12:0] Uout;
  input stop_i, start, start_cnt, clk, reset;
  output stop_o, st_out;
  wire   sw, start_temp, S2, n2, n57, n59, n61, n62, n63, n64, n65, n122, n123,
         n124, n126, n127, n128, n129, n130, n134, n136, n193, n194, n195,
         n197, n198, n199, n200, n201, n258, n259, n260, n262, n263, n264,
         n265, n266, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533;
  wire   [12:0] d1out;
  wire   [12:0] Q1;
  wire   [12:0] R1;
  wire   [12:0] r_mux;
  wire   [12:0] q_mux;
  wire   [12:0] U1;
  wire   [12:0] L1;
  wire   [12:0] l_mux;
  wire   [12:0] u_mux;
  wire   [12:0] d2out;
  wire   [12:0] d3out;
  wire   [12:0] d4out;
  wire   [12:0] R2;
  wire   [12:0] m1out;
  wire   [12:0] Q2;
  wire   [12:0] m2out;
  wire   [12:0] L2;
  wire   [12:0] m3out;
  wire   [12:0] U2;
  wire   [12:0] m4out;
  wire   [12:0] add1out;
  wire   [12:0] add2out;
  wire   [12:0] Q3;
  wire   [12:0] U3;

  DFFRHQX4 \Q2_reg[10]  ( .D(n330), .CK(clk), .RN(reset), .Q(Q2[10]) );
  DFFRHQX4 \R2_reg[12]  ( .D(n345), .CK(clk), .RN(reset), .Q(R2[12]) );
  degree_computation_1 degree1 ( .deg_Ri(deg_Ri), .deg_Qi(deg_Qi), .stop_i(
        stop_i), .d1out(d1out), .start(start), .deg_Ro(deg_Ro), .deg_Qo(deg_Qo), .stop_o(stop_o), .sw(sw), .clk(clk), .reset(reset) );
  mux_13_36 m1 ( .a(Q1), .b(R1), .sel(sw), .out(r_mux) );
  mux_13_35 m2 ( .a(R1), .b(Q1), .sel(sw), .out(q_mux) );
  mux_13_34 m3 ( .a(U1), .b(L1), .sel(sw), .out(l_mux) );
  mux_13_33 m4 ( .a(L1), .b(U1), .sel(sw), .out(u_mux) );
  feedback_ckt_7 D1 ( .Din(q_mux), .start(start_temp), .Qout(d1out), .clk(clk), 
        .reset(reset) );
  feedback_ckt_6 D2 ( .Din(r_mux), .start(start_temp), .Qout(d2out), .clk(clk), 
        .reset(reset) );
  feedback_ckt_5 D3 ( .Din(q_mux), .start(start_temp), .Qout(d3out), .clk(clk), 
        .reset(reset) );
  feedback_ckt_4 D4 ( .Din(r_mux), .start(n59), .Qout(d4out), .clk(clk), 
        .reset(reset) );
  multiplier_7 mx1 ( .a(R2), .b(d1out), .c(m1out) );
  multiplier_6 mx2 ( .a(d2out), .b(Q2), .c(m2out) );
  multiplier_5 mx3 ( .a(L2), .b(d3out), .c(m3out) );
  multiplier_4 mx4 ( .a(d4out), .b(U2), .c(m4out) );
  mux_13_32 m5 ( .a(R2), .b(add1out), .sel(n61), .out(Rout) );
  mux_13_31 m6 ( .a(Q2), .b(Q3), .sel(stop_i), .out(Qout) );
  mux_13_30 m7 ( .a(L2), .b(add2out), .sel(stop_i), .out(Lout) );
  mux_13_29 m8 ( .a(U2), .b(U3), .sel(n61), .out(Uout) );
  DFFRHQXL \R1_reg[12]  ( .D(n302), .CK(clk), .RN(reset), .Q(R1[12]) );
  DFFRHQXL \L1_reg[12]  ( .D(n359), .CK(clk), .RN(reset), .Q(L1[12]) );
  DFFRHQXL \R1_reg[2]  ( .D(n304), .CK(clk), .RN(reset), .Q(R1[2]) );
  DFFSX1 S3_reg ( .D(n416), .CK(clk), .SN(reset), .Q(st_out), .QN(n417) );
  DFFSX1 S2_reg ( .D(n301), .CK(clk), .SN(reset), .Q(S2) );
  DFFRHQX1 \Q3_reg[12]  ( .D(n346), .CK(clk), .RN(reset), .Q(Q3[12]) );
  DFFRHQX1 \Q3_reg[11]  ( .D(n347), .CK(clk), .RN(reset), .Q(Q3[11]) );
  DFFRHQX1 \Q3_reg[10]  ( .D(n348), .CK(clk), .RN(reset), .Q(Q3[10]) );
  DFFRHQX1 \Q3_reg[9]  ( .D(n349), .CK(clk), .RN(reset), .Q(Q3[9]) );
  DFFRHQX1 \Q3_reg[8]  ( .D(n350), .CK(clk), .RN(reset), .Q(Q3[8]) );
  DFFRHQX1 \Q3_reg[7]  ( .D(n351), .CK(clk), .RN(reset), .Q(Q3[7]) );
  DFFRHQX1 \Q3_reg[6]  ( .D(n352), .CK(clk), .RN(reset), .Q(Q3[6]) );
  DFFRHQX1 \Q3_reg[5]  ( .D(n353), .CK(clk), .RN(reset), .Q(Q3[5]) );
  DFFRHQX1 \Q3_reg[4]  ( .D(n354), .CK(clk), .RN(reset), .Q(Q3[4]) );
  DFFRHQX1 \Q3_reg[3]  ( .D(n355), .CK(clk), .RN(reset), .Q(Q3[3]) );
  DFFRHQX1 \Q3_reg[2]  ( .D(n356), .CK(clk), .RN(reset), .Q(Q3[2]) );
  DFFRHQX1 \Q3_reg[1]  ( .D(n357), .CK(clk), .RN(reset), .Q(Q3[1]) );
  DFFRHQX1 \Q3_reg[0]  ( .D(n358), .CK(clk), .RN(reset), .Q(Q3[0]) );
  DFFRHQX1 \U3_reg[12]  ( .D(n403), .CK(clk), .RN(reset), .Q(U3[12]) );
  DFFRHQX1 \U3_reg[11]  ( .D(n404), .CK(clk), .RN(reset), .Q(U3[11]) );
  DFFRHQX1 \U3_reg[10]  ( .D(n405), .CK(clk), .RN(reset), .Q(U3[10]) );
  DFFRHQX1 \U3_reg[9]  ( .D(n406), .CK(clk), .RN(reset), .Q(U3[9]) );
  DFFRHQX1 \U3_reg[8]  ( .D(n407), .CK(clk), .RN(reset), .Q(U3[8]) );
  DFFRHQX1 \U3_reg[7]  ( .D(n408), .CK(clk), .RN(reset), .Q(U3[7]) );
  DFFRHQX1 \U3_reg[6]  ( .D(n409), .CK(clk), .RN(reset), .Q(U3[6]) );
  DFFRHQX1 \U3_reg[5]  ( .D(n410), .CK(clk), .RN(reset), .Q(U3[5]) );
  DFFRHQX1 \U3_reg[4]  ( .D(n411), .CK(clk), .RN(reset), .Q(U3[4]) );
  DFFRHQX1 \U3_reg[3]  ( .D(n412), .CK(clk), .RN(reset), .Q(U3[3]) );
  DFFRHQX1 \U3_reg[2]  ( .D(n413), .CK(clk), .RN(reset), .Q(U3[2]) );
  DFFRHQX1 \U3_reg[1]  ( .D(n414), .CK(clk), .RN(reset), .Q(U3[1]) );
  DFFRHQX1 \U3_reg[0]  ( .D(n415), .CK(clk), .RN(reset), .Q(U3[0]) );
  DFFRHQX1 \R1_reg[1]  ( .D(n305), .CK(clk), .RN(reset), .Q(R1[1]) );
  DFFRHQX1 \R1_reg[0]  ( .D(n306), .CK(clk), .RN(reset), .Q(R1[0]) );
  DFFRHQX1 \Q1_reg[12]  ( .D(n307), .CK(clk), .RN(reset), .Q(Q1[12]) );
  DFFRHQX1 \Q1_reg[11]  ( .D(n308), .CK(clk), .RN(reset), .Q(Q1[11]) );
  DFFRHQX1 \Q1_reg[10]  ( .D(n309), .CK(clk), .RN(reset), .Q(Q1[10]) );
  DFFRHQX1 \Q1_reg[8]  ( .D(n311), .CK(clk), .RN(reset), .Q(Q1[8]) );
  DFFRHQX1 \Q1_reg[7]  ( .D(n312), .CK(clk), .RN(reset), .Q(Q1[7]) );
  DFFRHQX1 \Q1_reg[6]  ( .D(n313), .CK(clk), .RN(reset), .Q(Q1[6]) );
  DFFRHQX1 \Q1_reg[5]  ( .D(n314), .CK(clk), .RN(reset), .Q(Q1[5]) );
  DFFRHQX1 \Q1_reg[4]  ( .D(n315), .CK(clk), .RN(reset), .Q(Q1[4]) );
  DFFRHQX1 \Q1_reg[3]  ( .D(n316), .CK(clk), .RN(reset), .Q(Q1[3]) );
  DFFRHQX1 \Q1_reg[2]  ( .D(n317), .CK(clk), .RN(reset), .Q(Q1[2]) );
  DFFRHQX1 \Q1_reg[1]  ( .D(n318), .CK(clk), .RN(reset), .Q(Q1[1]) );
  DFFRHQX1 \Q1_reg[0]  ( .D(n319), .CK(clk), .RN(reset), .Q(Q1[0]) );
  DFFRHQX1 \L1_reg[2]  ( .D(n361), .CK(clk), .RN(reset), .Q(L1[2]) );
  DFFRHQX1 \L1_reg[1]  ( .D(n362), .CK(clk), .RN(reset), .Q(L1[1]) );
  DFFRHQX1 \L1_reg[0]  ( .D(n363), .CK(clk), .RN(reset), .Q(L1[0]) );
  DFFRHQX1 \U1_reg[12]  ( .D(n364), .CK(clk), .RN(reset), .Q(U1[12]) );
  DFFRHQX1 \U1_reg[11]  ( .D(n365), .CK(clk), .RN(reset), .Q(U1[11]) );
  DFFRHQX1 \U1_reg[10]  ( .D(n366), .CK(clk), .RN(reset), .Q(U1[10]) );
  DFFRHQX1 \U1_reg[8]  ( .D(n368), .CK(clk), .RN(reset), .Q(U1[8]) );
  DFFRHQX1 \U1_reg[7]  ( .D(n369), .CK(clk), .RN(reset), .Q(U1[7]) );
  DFFRHQX1 \U1_reg[6]  ( .D(n370), .CK(clk), .RN(reset), .Q(U1[6]) );
  DFFRHQX1 \U1_reg[5]  ( .D(n371), .CK(clk), .RN(reset), .Q(U1[5]) );
  DFFRHQX1 \U1_reg[4]  ( .D(n372), .CK(clk), .RN(reset), .Q(U1[4]) );
  DFFRHQX1 \U1_reg[3]  ( .D(n373), .CK(clk), .RN(reset), .Q(U1[3]) );
  DFFRHQX1 \U1_reg[2]  ( .D(n374), .CK(clk), .RN(reset), .Q(U1[2]) );
  DFFRHQX1 \U1_reg[1]  ( .D(n375), .CK(clk), .RN(reset), .Q(U1[1]) );
  DFFRHQX1 \U1_reg[0]  ( .D(n376), .CK(clk), .RN(reset), .Q(U1[0]) );
  DFFRHQX1 \Q1_reg[9]  ( .D(n310), .CK(clk), .RN(reset), .Q(Q1[9]) );
  DFFRHQX1 \U1_reg[9]  ( .D(n367), .CK(clk), .RN(reset), .Q(U1[9]) );
  DFFRHQX1 \R1_reg[7]  ( .D(n288), .CK(clk), .RN(reset), .Q(R1[7]) );
  DFFRHQX1 \R1_reg[4]  ( .D(n290), .CK(clk), .RN(reset), .Q(R1[4]) );
  DFFRHQX1 \L1_reg[5]  ( .D(n297), .CK(clk), .RN(reset), .Q(L1[5]) );
  DFFRHQX1 \L1_reg[4]  ( .D(n298), .CK(clk), .RN(reset), .Q(L1[4]) );
  DFFRHQX1 \R1_reg[9]  ( .D(n286), .CK(clk), .RN(reset), .Q(R1[9]) );
  DFFRHQX1 \L1_reg[9]  ( .D(n294), .CK(clk), .RN(reset), .Q(L1[9]) );
  DFFSX1 S1_reg ( .D(n300), .CK(clk), .SN(reset), .Q(start_temp), .QN(n2) );
  DFFRHQX1 \R2_reg[0]  ( .D(n333), .CK(clk), .RN(reset), .Q(R2[0]) );
  DFFRHQX1 \L2_reg[0]  ( .D(n390), .CK(clk), .RN(reset), .Q(L2[0]) );
  DFFRHQX1 \R2_reg[1]  ( .D(n334), .CK(clk), .RN(reset), .Q(R2[1]) );
  DFFRHQX1 \R2_reg[2]  ( .D(n335), .CK(clk), .RN(reset), .Q(R2[2]) );
  DFFRHQX1 \R2_reg[6]  ( .D(n339), .CK(clk), .RN(reset), .Q(R2[6]) );
  DFFRHQX1 \L2_reg[1]  ( .D(n391), .CK(clk), .RN(reset), .Q(L2[1]) );
  DFFRHQX1 \L2_reg[2]  ( .D(n392), .CK(clk), .RN(reset), .Q(L2[2]) );
  DFFRHQX1 \L2_reg[6]  ( .D(n396), .CK(clk), .RN(reset), .Q(L2[6]) );
  DFFRHQX1 \R2_reg[3]  ( .D(n336), .CK(clk), .RN(reset), .Q(R2[3]) );
  DFFRHQX1 \R2_reg[4]  ( .D(n337), .CK(clk), .RN(reset), .Q(R2[4]) );
  DFFRHQX1 \R2_reg[5]  ( .D(n338), .CK(clk), .RN(reset), .Q(R2[5]) );
  DFFRHQX1 \R2_reg[7]  ( .D(n340), .CK(clk), .RN(reset), .Q(R2[7]) );
  DFFRHQX1 \R2_reg[8]  ( .D(n341), .CK(clk), .RN(reset), .Q(R2[8]) );
  DFFRHQX1 \R2_reg[9]  ( .D(n342), .CK(clk), .RN(reset), .Q(R2[9]) );
  DFFRHQX1 \R2_reg[10]  ( .D(n343), .CK(clk), .RN(reset), .Q(R2[10]) );
  DFFRHQX1 \L2_reg[3]  ( .D(n393), .CK(clk), .RN(reset), .Q(L2[3]) );
  DFFRHQX1 \L2_reg[4]  ( .D(n394), .CK(clk), .RN(reset), .Q(L2[4]) );
  DFFRHQX1 \L2_reg[5]  ( .D(n395), .CK(clk), .RN(reset), .Q(L2[5]) );
  DFFRHQX1 \L2_reg[7]  ( .D(n397), .CK(clk), .RN(reset), .Q(L2[7]) );
  DFFRHQX1 \L2_reg[8]  ( .D(n398), .CK(clk), .RN(reset), .Q(L2[8]) );
  DFFRHQX1 \L2_reg[9]  ( .D(n399), .CK(clk), .RN(reset), .Q(L2[9]) );
  DFFRHQX1 \L2_reg[10]  ( .D(n400), .CK(clk), .RN(reset), .Q(L2[10]) );
  DFFRHQX1 \Q2_reg[2]  ( .D(n322), .CK(clk), .RN(reset), .Q(Q2[2]) );
  DFFRHQX1 \Q2_reg[6]  ( .D(n326), .CK(clk), .RN(reset), .Q(Q2[6]) );
  DFFRHQX1 \Q2_reg[8]  ( .D(n328), .CK(clk), .RN(reset), .Q(Q2[8]) );
  DFFRHQX1 \Q2_reg[12]  ( .D(n332), .CK(clk), .RN(reset), .Q(Q2[12]) );
  DFFRHQX1 \U2_reg[2]  ( .D(n379), .CK(clk), .RN(reset), .Q(U2[2]) );
  DFFRHQX1 \U2_reg[5]  ( .D(n382), .CK(clk), .RN(reset), .Q(U2[5]) );
  DFFRHQX1 \U2_reg[6]  ( .D(n383), .CK(clk), .RN(reset), .Q(U2[6]) );
  DFFRHQX1 \U2_reg[7]  ( .D(n384), .CK(clk), .RN(reset), .Q(U2[7]) );
  DFFRHQX1 \U2_reg[8]  ( .D(n385), .CK(clk), .RN(reset), .Q(U2[8]) );
  DFFRHQX1 \U2_reg[12]  ( .D(n389), .CK(clk), .RN(reset), .Q(U2[12]) );
  DFFRHQX1 \Q2_reg[9]  ( .D(n329), .CK(clk), .RN(reset), .Q(Q2[9]) );
  DFFRHQX1 \U2_reg[9]  ( .D(n386), .CK(clk), .RN(reset), .Q(U2[9]) );
  DFFRHQX1 \Q2_reg[0]  ( .D(n320), .CK(clk), .RN(reset), .Q(Q2[0]) );
  DFFRHQX1 \U2_reg[0]  ( .D(n377), .CK(clk), .RN(reset), .Q(U2[0]) );
  DFFRHQX1 \Q2_reg[1]  ( .D(n321), .CK(clk), .RN(reset), .Q(Q2[1]) );
  DFFRHQX1 \U2_reg[1]  ( .D(n378), .CK(clk), .RN(reset), .Q(U2[1]) );
  DFFRHQXL \R1_reg[11]  ( .D(n284), .CK(clk), .RN(reset), .Q(R1[11]) );
  DFFRHQXL \R1_reg[10]  ( .D(n285), .CK(clk), .RN(reset), .Q(R1[10]) );
  DFFRHQXL \R1_reg[8]  ( .D(n287), .CK(clk), .RN(reset), .Q(R1[8]) );
  DFFRHQXL \R1_reg[3]  ( .D(n291), .CK(clk), .RN(reset), .Q(R1[3]) );
  DFFRHQXL \L1_reg[11]  ( .D(n292), .CK(clk), .RN(reset), .Q(L1[11]) );
  DFFRHQXL \L1_reg[10]  ( .D(n293), .CK(clk), .RN(reset), .Q(L1[10]) );
  DFFRHQXL \L1_reg[8]  ( .D(n295), .CK(clk), .RN(reset), .Q(L1[8]) );
  DFFRHQXL \L1_reg[7]  ( .D(n296), .CK(clk), .RN(reset), .Q(L1[7]) );
  DFFRHQXL \L1_reg[3]  ( .D(n299), .CK(clk), .RN(reset), .Q(L1[3]) );
  DFFRHQX2 \Q2_reg[11]  ( .D(n331), .CK(clk), .RN(reset), .Q(Q2[11]) );
  DFFRHQXL \R1_reg[5]  ( .D(n289), .CK(clk), .RN(reset), .Q(R1[5]) );
  DFFRHQX2 \L2_reg[11]  ( .D(n401), .CK(clk), .RN(reset), .Q(L2[11]) );
  DFFRHQXL \R1_reg[6]  ( .D(n303), .CK(clk), .RN(reset), .Q(R1[6]) );
  DFFRHQX2 \Q2_reg[4]  ( .D(n324), .CK(clk), .RN(reset), .Q(Q2[4]) );
  DFFRHQX2 \U2_reg[10]  ( .D(n387), .CK(clk), .RN(reset), .Q(U2[10]) );
  DFFRHQX2 \U2_reg[3]  ( .D(n380), .CK(clk), .RN(reset), .Q(U2[3]) );
  DFFRHQX2 \Q2_reg[3]  ( .D(n323), .CK(clk), .RN(reset), .Q(Q2[3]) );
  DFFRHQX2 \U2_reg[11]  ( .D(n388), .CK(clk), .RN(reset), .Q(U2[11]) );
  DFFRHQX2 \L2_reg[12]  ( .D(n402), .CK(clk), .RN(reset), .Q(L2[12]) );
  DFFRHQX2 \U2_reg[4]  ( .D(n381), .CK(clk), .RN(reset), .Q(U2[4]) );
  DFFRHQX2 \R2_reg[11]  ( .D(n344), .CK(clk), .RN(reset), .Q(R2[11]) );
  DFFRHQXL \L1_reg[6]  ( .D(n360), .CK(clk), .RN(reset), .Q(L1[6]) );
  DFFRHQX2 \Q2_reg[5]  ( .D(n325), .CK(clk), .RN(reset), .Q(Q2[5]) );
  DFFRHQX2 \Q2_reg[7]  ( .D(n327), .CK(clk), .RN(reset), .Q(Q2[7]) );
  MX2X2 U2_inst ( .A(Rin[5]), .B(R1[5]), .S0(n199), .Y(n289) );
  INVX1 U3_inst ( .A(R1[12]), .Y(n57) );
  AOI2BB2X1 U4 ( .B0(Rin[12]), .B1(n262), .A0N(n57), .A1N(n275), .Y(n420) );
  MX2X1 U5 ( .A(L1[5]), .B(Lin[5]), .S0(n65), .Y(n297) );
  MX2X1 U6 ( .A(R1[4]), .B(Rin[4]), .S0(n65), .Y(n290) );
  MX2X1 U7 ( .A(R1[7]), .B(Rin[7]), .S0(n275), .Y(n288) );
  XOR2X1 U8 ( .A(m4out[8]), .B(m3out[8]), .Y(add2out[8]) );
  XOR2X1 U9 ( .A(m4out[11]), .B(m3out[11]), .Y(add2out[11]) );
  XOR2X1 U10 ( .A(m2out[5]), .B(m1out[5]), .Y(add1out[5]) );
  XOR2X1 U11 ( .A(m4out[5]), .B(m3out[5]), .Y(add2out[5]) );
  MX2X1 U12 ( .A(L1[8]), .B(Lin[8]), .S0(n65), .Y(n295) );
  MX2X1 U13 ( .A(L1[7]), .B(Lin[7]), .S0(n65), .Y(n296) );
  MX2X1 U14 ( .A(L1[10]), .B(Lin[10]), .S0(n65), .Y(n293) );
  MX2X1 U15 ( .A(L1[3]), .B(Lin[3]), .S0(n65), .Y(n299) );
  MX2X1 U16 ( .A(R1[3]), .B(Rin[3]), .S0(n65), .Y(n291) );
  MX2X1 U17 ( .A(L1[4]), .B(Lin[4]), .S0(n65), .Y(n298) );
  MX2X1 U18 ( .A(L1[11]), .B(Lin[11]), .S0(n65), .Y(n292) );
  MX2X1 U19 ( .A(R1[8]), .B(Rin[8]), .S0(n277), .Y(n287) );
  MX2X1 U20 ( .A(R1[10]), .B(Rin[10]), .S0(n276), .Y(n285) );
  MX2X1 U21 ( .A(R1[11]), .B(Rin[11]), .S0(n260), .Y(n284) );
  MX2X1 U22 ( .A(R1[9]), .B(Rin[9]), .S0(n271), .Y(n286) );
  INVXL U23 ( .A(n420), .Y(n302) );
  INVXL U24 ( .A(n477), .Y(n359) );
  INVXL U25 ( .A(n422), .Y(n304) );
  INVXL U26 ( .A(n423), .Y(n305) );
  INVXL U27 ( .A(n421), .Y(n303) );
  INVXL U28 ( .A(n479), .Y(n361) );
  INVXL U29 ( .A(n480), .Y(n362) );
  INVXL U30 ( .A(n478), .Y(n360) );
  AOI22XL U31 ( .A0(n195), .A1(U2[12]), .B0(u_mux[12]), .B1(n262), .Y(n507) );
  AOI22XL U32 ( .A0(n199), .A1(U2[9]), .B0(u_mux[9]), .B1(n275), .Y(n504) );
  AOI22XL U33 ( .A0(n194), .A1(U2[8]), .B0(u_mux[8]), .B1(n274), .Y(n503) );
  AOI22XL U34 ( .A0(n199), .A1(U2[7]), .B0(u_mux[7]), .B1(n271), .Y(n502) );
  AOI22XL U35 ( .A0(n198), .A1(U2[6]), .B0(u_mux[6]), .B1(n271), .Y(n501) );
  AOI22XL U36 ( .A0(n198), .A1(U2[5]), .B0(u_mux[5]), .B1(n259), .Y(n500) );
  AOI22XL U37 ( .A0(n136), .A1(U2[4]), .B0(u_mux[4]), .B1(n266), .Y(n499) );
  AOI22XL U38 ( .A0(n195), .A1(U2[1]), .B0(u_mux[1]), .B1(n266), .Y(n496) );
  AOI22XL U39 ( .A0(n193), .A1(U2[0]), .B0(u_mux[0]), .B1(n265), .Y(n495) );
  AOI22XL U40 ( .A0(R2[10]), .A1(n123), .B0(r_mux[10]), .B1(n277), .Y(n461) );
  AOI22XL U41 ( .A0(R2[9]), .A1(n127), .B0(r_mux[9]), .B1(n270), .Y(n460) );
  AOI22XL U42 ( .A0(R2[8]), .A1(n124), .B0(r_mux[8]), .B1(n262), .Y(n459) );
  AOI22XL U43 ( .A0(R2[7]), .A1(n200), .B0(r_mux[7]), .B1(n271), .Y(n458) );
  AOI22XL U44 ( .A0(R2[6]), .A1(n198), .B0(r_mux[6]), .B1(n260), .Y(n457) );
  AOI22XL U45 ( .A0(R2[5]), .A1(n258), .B0(r_mux[5]), .B1(n259), .Y(n456) );
  AOI22XL U46 ( .A0(R2[4]), .A1(n199), .B0(r_mux[4]), .B1(n274), .Y(n455) );
  AOI22XL U47 ( .A0(R2[3]), .A1(n124), .B0(r_mux[3]), .B1(n259), .Y(n454) );
  AOI22XL U48 ( .A0(n130), .A1(Q2[12]), .B0(q_mux[12]), .B1(n260), .Y(n450) );
  AOI22XL U49 ( .A0(n130), .A1(Q2[9]), .B0(q_mux[9]), .B1(n260), .Y(n447) );
  AOI22XL U50 ( .A0(n134), .A1(Q2[8]), .B0(q_mux[8]), .B1(n262), .Y(n446) );
  AOI22XL U51 ( .A0(n130), .A1(Q2[7]), .B0(q_mux[7]), .B1(n263), .Y(n445) );
  AOI22XL U52 ( .A0(n129), .A1(Q2[6]), .B0(q_mux[6]), .B1(n260), .Y(n444) );
  AOI22XL U53 ( .A0(n127), .A1(Q2[5]), .B0(q_mux[5]), .B1(n260), .Y(n443) );
  AOI22XL U54 ( .A0(n129), .A1(Q2[4]), .B0(q_mux[4]), .B1(n259), .Y(n442) );
  AOI22XL U55 ( .A0(n128), .A1(Q2[1]), .B0(q_mux[1]), .B1(n264), .Y(n439) );
  AOI22XL U56 ( .A0(n129), .A1(Q2[0]), .B0(q_mux[0]), .B1(n263), .Y(n438) );
  AOI22XL U57 ( .A0(n275), .A1(Q2[1]), .B0(Q3[1]), .B1(n201), .Y(n475) );
  AOI22XL U58 ( .A0(L2[12]), .A1(n201), .B0(l_mux[12]), .B1(n264), .Y(n520) );
  AOI22XL U59 ( .A0(n200), .A1(U2[11]), .B0(u_mux[11]), .B1(n265), .Y(n506) );
  AOI22XL U60 ( .A0(n193), .A1(U2[10]), .B0(u_mux[10]), .B1(n271), .Y(n505) );
  AOI22XL U61 ( .A0(n197), .A1(U2[3]), .B0(u_mux[3]), .B1(n272), .Y(n498) );
  AOI22XL U62 ( .A0(R2[12]), .A1(n193), .B0(r_mux[12]), .B1(n273), .Y(n463) );
  AOI22XL U63 ( .A0(R2[11]), .A1(n127), .B0(r_mux[11]), .B1(n272), .Y(n462) );
  AOI22XL U64 ( .A0(n130), .A1(Q2[11]), .B0(q_mux[11]), .B1(n260), .Y(n449) );
  AOI22XL U65 ( .A0(n136), .A1(Q2[10]), .B0(q_mux[10]), .B1(n275), .Y(n448) );
  AOI22XL U66 ( .A0(n128), .A1(Q2[3]), .B0(q_mux[3]), .B1(n262), .Y(n441) );
  AOI22XL U67 ( .A0(n273), .A1(U2[0]), .B0(U3[0]), .B1(n201), .Y(n533) );
  AOI22XL U68 ( .A0(n272), .A1(U2[1]), .B0(U3[1]), .B1(n258), .Y(n532) );
  AOI22XL U69 ( .A0(L2[9]), .A1(n199), .B0(l_mux[9]), .B1(n274), .Y(n517) );
  AOI22XL U70 ( .A0(L2[8]), .A1(n197), .B0(l_mux[8]), .B1(n273), .Y(n516) );
  AOI22XL U71 ( .A0(L2[5]), .A1(n123), .B0(l_mux[5]), .B1(n262), .Y(n513) );
  AOI22XL U72 ( .A0(L2[3]), .A1(n200), .B0(l_mux[3]), .B1(n275), .Y(n511) );
  AOI22XL U73 ( .A0(n274), .A1(U2[3]), .B0(U3[3]), .B1(n280), .Y(n530) );
  AOI22XL U74 ( .A0(n63), .A1(U2[4]), .B0(U3[4]), .B1(n201), .Y(n529) );
  AOI22XL U75 ( .A0(n266), .A1(U2[5]), .B0(U3[5]), .B1(n201), .Y(n528) );
  AOI22XL U76 ( .A0(n272), .A1(U2[6]), .B0(U3[6]), .B1(n258), .Y(n527) );
  AOI22XL U77 ( .A0(n259), .A1(U2[7]), .B0(U3[7]), .B1(n258), .Y(n526) );
  AOI22XL U78 ( .A0(n264), .A1(U2[8]), .B0(U3[8]), .B1(n258), .Y(n525) );
  AOI22XL U79 ( .A0(n277), .A1(U2[9]), .B0(U3[9]), .B1(n258), .Y(n524) );
  AOI22XL U80 ( .A0(n260), .A1(U2[10]), .B0(U3[10]), .B1(n258), .Y(n523) );
  AOI22XL U81 ( .A0(n270), .A1(U2[11]), .B0(U3[11]), .B1(n201), .Y(n522) );
  AOI22XL U82 ( .A0(n276), .A1(U2[12]), .B0(U3[12]), .B1(n278), .Y(n521) );
  AOI22XL U83 ( .A0(n272), .A1(Q2[0]), .B0(Q3[0]), .B1(n201), .Y(n476) );
  AOI22XL U84 ( .A0(n275), .A1(Q2[3]), .B0(Q3[3]), .B1(n278), .Y(n473) );
  AOI22XL U85 ( .A0(n273), .A1(Q2[4]), .B0(Q3[4]), .B1(n280), .Y(n472) );
  AOI22XL U86 ( .A0(n63), .A1(Q2[5]), .B0(Q3[5]), .B1(n200), .Y(n471) );
  AOI22XL U87 ( .A0(n259), .A1(Q2[6]), .B0(Q3[6]), .B1(n281), .Y(n470) );
  AOI22XL U88 ( .A0(n271), .A1(Q2[9]), .B0(Q3[9]), .B1(n278), .Y(n467) );
  AOI22XL U89 ( .A0(n265), .A1(Q2[12]), .B0(Q3[12]), .B1(n279), .Y(n464) );
  AOI22XL U90 ( .A0(n265), .A1(Q2[7]), .B0(Q3[7]), .B1(n279), .Y(n469) );
  AOI22XL U91 ( .A0(n260), .A1(Q2[8]), .B0(Q3[8]), .B1(n279), .Y(n468) );
  AOI22XL U92 ( .A0(n270), .A1(Q2[10]), .B0(Q3[10]), .B1(n279), .Y(n466) );
  AOI22XL U93 ( .A0(n274), .A1(Q2[11]), .B0(Q3[11]), .B1(n278), .Y(n465) );
  AOI22XL U94 ( .A0(L2[11]), .A1(n122), .B0(l_mux[11]), .B1(n263), .Y(n519) );
  AOI22XL U95 ( .A0(L2[10]), .A1(n258), .B0(l_mux[10]), .B1(n276), .Y(n518) );
  INVX1 U96 ( .A(n64), .Y(n65) );
  INVX1 U97 ( .A(n270), .Y(n126) );
  INVX1 U98 ( .A(n266), .Y(n127) );
  INVX1 U99 ( .A(n273), .Y(n124) );
  INVX1 U100 ( .A(n274), .Y(n123) );
  INVX1 U101 ( .A(n274), .Y(n122) );
  INVX1 U102 ( .A(n262), .Y(n199) );
  INVX1 U103 ( .A(n262), .Y(n198) );
  INVX1 U104 ( .A(n263), .Y(n197) );
  INVX1 U105 ( .A(n263), .Y(n195) );
  INVX1 U106 ( .A(n264), .Y(n193) );
  INVX1 U107 ( .A(n264), .Y(n136) );
  INVX1 U108 ( .A(n265), .Y(n130) );
  INVX1 U109 ( .A(n265), .Y(n129) );
  INVX1 U110 ( .A(n264), .Y(n134) );
  INVX1 U111 ( .A(n266), .Y(n128) );
  INVX1 U112 ( .A(n263), .Y(n194) );
  INVX1 U113 ( .A(n262), .Y(n200) );
  INVX1 U114 ( .A(n259), .Y(n258) );
  INVX1 U115 ( .A(n260), .Y(n201) );
  INVX1 U116 ( .A(n281), .Y(n259) );
  INVX1 U117 ( .A(n279), .Y(n270) );
  INVX1 U118 ( .A(n280), .Y(n262) );
  INVX1 U119 ( .A(n281), .Y(n260) );
  INVX1 U120 ( .A(n281), .Y(n274) );
  INVX1 U121 ( .A(n278), .Y(n271) );
  INVX1 U122 ( .A(n280), .Y(n273) );
  INVX1 U123 ( .A(n279), .Y(n272) );
  INVX1 U124 ( .A(n279), .Y(n275) );
  INVX1 U125 ( .A(n280), .Y(n264) );
  INVX1 U126 ( .A(n279), .Y(n266) );
  INVX1 U127 ( .A(n279), .Y(n265) );
  INVX1 U128 ( .A(n278), .Y(n276) );
  INVX1 U129 ( .A(n278), .Y(n277) );
  INVX1 U130 ( .A(n280), .Y(n263) );
  INVX1 U131 ( .A(n63), .Y(n281) );
  INVX1 U132 ( .A(n63), .Y(n279) );
  INVX1 U133 ( .A(n63), .Y(n278) );
  INVX1 U134 ( .A(n63), .Y(n280) );
  INVX1 U135 ( .A(n64), .Y(n63) );
  INVX1 U136 ( .A(start_cnt), .Y(n64) );
  XOR2X1 U137 ( .A(m3out[10]), .B(m4out[10]), .Y(add2out[10]) );
  XOR2X1 U138 ( .A(m1out[10]), .B(m2out[10]), .Y(add1out[10]) );
  XOR2X1 U139 ( .A(m1out[8]), .B(m2out[8]), .Y(add1out[8]) );
  XOR2X1 U140 ( .A(m1out[4]), .B(m2out[4]), .Y(add1out[4]) );
  XOR2X1 U141 ( .A(m4out[6]), .B(m3out[6]), .Y(add2out[6]) );
  XOR2X1 U142 ( .A(m2out[6]), .B(m1out[6]), .Y(add1out[6]) );
  XOR2X1 U143 ( .A(m4out[2]), .B(m3out[2]), .Y(add2out[2]) );
  XOR2X1 U144 ( .A(m4out[1]), .B(m3out[1]), .Y(add2out[1]) );
  XOR2X1 U145 ( .A(m2out[1]), .B(m1out[1]), .Y(add1out[1]) );
  XOR2X1 U146 ( .A(m2out[2]), .B(m1out[2]), .Y(add1out[2]) );
  XOR2X1 U147 ( .A(m2out[12]), .B(m1out[12]), .Y(add1out[12]) );
  XOR2X1 U148 ( .A(m4out[12]), .B(m3out[12]), .Y(add2out[12]) );
  XOR2X1 U149 ( .A(m1out[7]), .B(m2out[7]), .Y(add1out[7]) );
  XOR2X1 U150 ( .A(m3out[7]), .B(m4out[7]), .Y(add2out[7]) );
  XOR2X1 U151 ( .A(m3out[3]), .B(m4out[3]), .Y(add2out[3]) );
  XOR2X1 U152 ( .A(m3out[4]), .B(m4out[4]), .Y(add2out[4]) );
  XOR2X1 U153 ( .A(m3out[9]), .B(m4out[9]), .Y(add2out[9]) );
  XOR2X1 U154 ( .A(m1out[3]), .B(m2out[3]), .Y(add1out[3]) );
  XOR2X1 U155 ( .A(m1out[9]), .B(m2out[9]), .Y(add1out[9]) );
  XOR2X1 U156 ( .A(m1out[11]), .B(m2out[11]), .Y(add1out[11]) );
  XOR2X1 U157 ( .A(m2out[0]), .B(m1out[0]), .Y(add1out[0]) );
  XOR2X1 U158 ( .A(m4out[0]), .B(m3out[0]), .Y(add2out[0]) );
  INVX1 U159 ( .A(n2), .Y(n59) );
  INVX1 U160 ( .A(n62), .Y(n61) );
  INVX1 U161 ( .A(n520), .Y(n402) );
  INVX1 U162 ( .A(n518), .Y(n400) );
  MXI2X1 U163 ( .A(n283), .B(n282), .S0(n65), .Y(n294) );
  INVX1 U164 ( .A(L1[9]), .Y(n283) );
  INVX1 U165 ( .A(Lin[9]), .Y(n282) );
  OAI2BB2X1 U166 ( .B0(n63), .B1(n417), .A0N(S2), .A1N(n276), .Y(n416) );
  AOI22X1 U167 ( .A0(R1[2]), .A1(n122), .B0(Rin[2]), .B1(n265), .Y(n422) );
  AOI22X1 U168 ( .A0(L1[12]), .A1(n129), .B0(Lin[12]), .B1(n264), .Y(n477) );
  INVX1 U169 ( .A(n519), .Y(n401) );
  INVX1 U170 ( .A(n532), .Y(n414) );
  INVX1 U171 ( .A(n496), .Y(n378) );
  INVX1 U172 ( .A(n475), .Y(n357) );
  INVX1 U173 ( .A(n439), .Y(n321) );
  INVX1 U174 ( .A(n533), .Y(n415) );
  INVX1 U175 ( .A(n495), .Y(n377) );
  INVX1 U176 ( .A(n476), .Y(n358) );
  INVX1 U177 ( .A(n438), .Y(n320) );
  INVX1 U178 ( .A(n524), .Y(n406) );
  INVX1 U179 ( .A(n504), .Y(n386) );
  INVX1 U180 ( .A(n467), .Y(n349) );
  INVX1 U181 ( .A(n447), .Y(n329) );
  INVX1 U182 ( .A(n531), .Y(n413) );
  AOI22X1 U183 ( .A0(n262), .A1(U2[2]), .B0(U3[2]), .B1(n258), .Y(n531) );
  INVX1 U184 ( .A(n530), .Y(n412) );
  INVX1 U185 ( .A(n529), .Y(n411) );
  INVX1 U186 ( .A(n528), .Y(n410) );
  INVX1 U187 ( .A(n527), .Y(n409) );
  INVX1 U188 ( .A(n526), .Y(n408) );
  INVX1 U189 ( .A(n525), .Y(n407) );
  INVX1 U190 ( .A(n523), .Y(n405) );
  INVX1 U191 ( .A(n522), .Y(n404) );
  INVX1 U192 ( .A(n521), .Y(n403) );
  INVX1 U193 ( .A(n507), .Y(n389) );
  INVX1 U194 ( .A(n506), .Y(n388) );
  INVX1 U195 ( .A(n505), .Y(n387) );
  INVX1 U196 ( .A(n503), .Y(n385) );
  INVX1 U197 ( .A(n502), .Y(n384) );
  INVX1 U198 ( .A(n501), .Y(n383) );
  INVX1 U199 ( .A(n500), .Y(n382) );
  INVX1 U200 ( .A(n499), .Y(n381) );
  INVX1 U201 ( .A(n498), .Y(n380) );
  INVX1 U202 ( .A(n497), .Y(n379) );
  AOI22X1 U203 ( .A0(n197), .A1(U2[2]), .B0(u_mux[2]), .B1(n270), .Y(n497) );
  INVX1 U204 ( .A(n474), .Y(n356) );
  AOI22X1 U205 ( .A0(n263), .A1(Q2[2]), .B0(Q3[2]), .B1(n278), .Y(n474) );
  INVX1 U206 ( .A(n473), .Y(n355) );
  INVX1 U207 ( .A(n472), .Y(n354) );
  INVX1 U208 ( .A(n471), .Y(n353) );
  INVX1 U209 ( .A(n470), .Y(n352) );
  INVX1 U210 ( .A(n469), .Y(n351) );
  INVX1 U211 ( .A(n468), .Y(n350) );
  INVX1 U212 ( .A(n466), .Y(n348) );
  INVX1 U213 ( .A(n465), .Y(n347) );
  INVX1 U214 ( .A(n464), .Y(n346) );
  INVX1 U215 ( .A(n450), .Y(n332) );
  INVX1 U216 ( .A(n449), .Y(n331) );
  INVX1 U217 ( .A(n448), .Y(n330) );
  INVX1 U218 ( .A(n446), .Y(n328) );
  INVX1 U219 ( .A(n445), .Y(n327) );
  INVX1 U220 ( .A(n444), .Y(n326) );
  INVX1 U221 ( .A(n443), .Y(n325) );
  INVX1 U222 ( .A(n442), .Y(n324) );
  INVX1 U223 ( .A(n441), .Y(n323) );
  INVX1 U224 ( .A(n440), .Y(n322) );
  AOI22X1 U225 ( .A0(n134), .A1(Q2[2]), .B0(q_mux[2]), .B1(n276), .Y(n440) );
  INVX1 U226 ( .A(n517), .Y(n399) );
  INVX1 U227 ( .A(n516), .Y(n398) );
  INVX1 U228 ( .A(n515), .Y(n397) );
  AOI22X1 U229 ( .A0(L2[7]), .A1(n123), .B0(l_mux[7]), .B1(n277), .Y(n515) );
  INVX1 U230 ( .A(n514), .Y(n396) );
  AOI22X1 U231 ( .A0(L2[6]), .A1(n128), .B0(l_mux[6]), .B1(n272), .Y(n514) );
  INVX1 U232 ( .A(n513), .Y(n395) );
  INVX1 U233 ( .A(n512), .Y(n394) );
  AOI22X1 U234 ( .A0(L2[4]), .A1(n134), .B0(l_mux[4]), .B1(n272), .Y(n512) );
  INVX1 U235 ( .A(n511), .Y(n393) );
  INVX1 U236 ( .A(n510), .Y(n392) );
  AOI22X1 U237 ( .A0(L2[2]), .A1(n124), .B0(l_mux[2]), .B1(n276), .Y(n510) );
  INVX1 U238 ( .A(n509), .Y(n391) );
  AOI22X1 U239 ( .A0(L2[1]), .A1(n128), .B0(l_mux[1]), .B1(n266), .Y(n509) );
  INVX1 U240 ( .A(n508), .Y(n390) );
  AOI22X1 U241 ( .A0(L2[0]), .A1(n194), .B0(l_mux[0]), .B1(n265), .Y(n508) );
  INVX1 U242 ( .A(n494), .Y(n376) );
  AOI22X1 U243 ( .A0(U1[0]), .A1(n198), .B0(Uin[0]), .B1(n276), .Y(n494) );
  INVX1 U244 ( .A(n493), .Y(n375) );
  AOI22X1 U245 ( .A0(U1[1]), .A1(n124), .B0(Uin[1]), .B1(n271), .Y(n493) );
  INVX1 U246 ( .A(n492), .Y(n374) );
  AOI22X1 U247 ( .A0(U1[2]), .A1(n129), .B0(Uin[2]), .B1(n270), .Y(n492) );
  INVX1 U248 ( .A(n491), .Y(n373) );
  AOI22X1 U249 ( .A0(U1[3]), .A1(n124), .B0(Uin[3]), .B1(n276), .Y(n491) );
  INVX1 U250 ( .A(n490), .Y(n372) );
  AOI22X1 U251 ( .A0(U1[4]), .A1(n134), .B0(Uin[4]), .B1(n270), .Y(n490) );
  INVX1 U252 ( .A(n489), .Y(n371) );
  AOI22X1 U253 ( .A0(U1[5]), .A1(n193), .B0(Uin[5]), .B1(n277), .Y(n489) );
  INVX1 U254 ( .A(n488), .Y(n370) );
  AOI22X1 U255 ( .A0(U1[6]), .A1(n126), .B0(Uin[6]), .B1(n273), .Y(n488) );
  INVX1 U256 ( .A(n487), .Y(n369) );
  AOI22X1 U257 ( .A0(U1[7]), .A1(n194), .B0(Uin[7]), .B1(n275), .Y(n487) );
  INVX1 U258 ( .A(n486), .Y(n368) );
  AOI22X1 U259 ( .A0(U1[8]), .A1(n126), .B0(Uin[8]), .B1(n274), .Y(n486) );
  INVX1 U260 ( .A(n485), .Y(n367) );
  AOI22X1 U261 ( .A0(U1[9]), .A1(n195), .B0(Uin[9]), .B1(n264), .Y(n485) );
  INVX1 U262 ( .A(n484), .Y(n366) );
  AOI22X1 U263 ( .A0(U1[10]), .A1(n194), .B0(Uin[10]), .B1(n273), .Y(n484) );
  INVX1 U264 ( .A(n483), .Y(n365) );
  AOI22X1 U265 ( .A0(U1[11]), .A1(n197), .B0(Uin[11]), .B1(n274), .Y(n483) );
  INVX1 U266 ( .A(n482), .Y(n364) );
  AOI22X1 U267 ( .A0(U1[12]), .A1(n126), .B0(Uin[12]), .B1(n275), .Y(n482) );
  INVX1 U268 ( .A(n481), .Y(n363) );
  AOI22X1 U269 ( .A0(L1[0]), .A1(n130), .B0(Lin[0]), .B1(n273), .Y(n481) );
  AOI22X1 U270 ( .A0(L1[1]), .A1(n126), .B0(Lin[1]), .B1(n263), .Y(n480) );
  INVX1 U271 ( .A(n463), .Y(n345) );
  INVX1 U272 ( .A(n462), .Y(n344) );
  INVX1 U273 ( .A(n461), .Y(n343) );
  INVX1 U274 ( .A(n460), .Y(n342) );
  INVX1 U275 ( .A(n459), .Y(n341) );
  INVX1 U276 ( .A(n458), .Y(n340) );
  INVX1 U277 ( .A(n457), .Y(n339) );
  INVX1 U278 ( .A(n456), .Y(n338) );
  INVX1 U279 ( .A(n455), .Y(n337) );
  INVX1 U280 ( .A(n454), .Y(n336) );
  INVX1 U281 ( .A(n453), .Y(n335) );
  AOI22X1 U282 ( .A0(R2[2]), .A1(n124), .B0(r_mux[2]), .B1(n277), .Y(n453) );
  INVX1 U283 ( .A(n452), .Y(n334) );
  AOI22X1 U284 ( .A0(R2[1]), .A1(n195), .B0(r_mux[1]), .B1(n63), .Y(n452) );
  INVX1 U285 ( .A(n451), .Y(n333) );
  AOI22X1 U286 ( .A0(R2[0]), .A1(n122), .B0(r_mux[0]), .B1(n263), .Y(n451) );
  INVX1 U287 ( .A(n437), .Y(n319) );
  AOI22X1 U288 ( .A0(Q1[0]), .A1(n195), .B0(Qin[0]), .B1(n274), .Y(n437) );
  INVX1 U289 ( .A(n436), .Y(n318) );
  AOI22X1 U290 ( .A0(Q1[1]), .A1(n136), .B0(Qin[1]), .B1(n272), .Y(n436) );
  INVX1 U291 ( .A(n435), .Y(n317) );
  AOI22X1 U292 ( .A0(Q1[2]), .A1(n127), .B0(Qin[2]), .B1(n270), .Y(n435) );
  INVX1 U293 ( .A(n434), .Y(n316) );
  AOI22X1 U294 ( .A0(Q1[3]), .A1(n193), .B0(Qin[3]), .B1(n271), .Y(n434) );
  INVX1 U295 ( .A(n433), .Y(n315) );
  AOI22X1 U296 ( .A0(Q1[4]), .A1(n258), .B0(Qin[4]), .B1(n277), .Y(n433) );
  INVX1 U297 ( .A(n432), .Y(n314) );
  AOI22X1 U298 ( .A0(Q1[5]), .A1(n124), .B0(Qin[5]), .B1(n276), .Y(n432) );
  INVX1 U299 ( .A(n431), .Y(n313) );
  AOI22X1 U300 ( .A0(Q1[6]), .A1(n123), .B0(Qin[6]), .B1(n264), .Y(n431) );
  INVX1 U301 ( .A(n430), .Y(n312) );
  AOI22X1 U302 ( .A0(Q1[7]), .A1(n122), .B0(Qin[7]), .B1(n271), .Y(n430) );
  INVX1 U303 ( .A(n429), .Y(n311) );
  AOI22X1 U304 ( .A0(Q1[8]), .A1(n278), .B0(Qin[8]), .B1(n266), .Y(n429) );
  INVX1 U305 ( .A(n428), .Y(n310) );
  AOI22X1 U306 ( .A0(Q1[9]), .A1(n278), .B0(Qin[9]), .B1(n259), .Y(n428) );
  INVX1 U307 ( .A(n427), .Y(n309) );
  AOI22X1 U308 ( .A0(Q1[10]), .A1(n123), .B0(Qin[10]), .B1(n275), .Y(n427) );
  INVX1 U309 ( .A(n426), .Y(n308) );
  AOI22X1 U310 ( .A0(Q1[11]), .A1(n122), .B0(Qin[11]), .B1(n263), .Y(n426) );
  INVX1 U311 ( .A(n425), .Y(n307) );
  AOI22X1 U312 ( .A0(Q1[12]), .A1(n123), .B0(Qin[12]), .B1(n266), .Y(n425) );
  INVX1 U313 ( .A(n424), .Y(n306) );
  AOI22X1 U314 ( .A0(R1[0]), .A1(n123), .B0(Rin[0]), .B1(n265), .Y(n424) );
  AOI22X1 U315 ( .A0(R1[1]), .A1(n122), .B0(Rin[1]), .B1(n264), .Y(n423) );
  AOI22X1 U316 ( .A0(L1[6]), .A1(n134), .B0(Lin[6]), .B1(n272), .Y(n478) );
  AOI22X1 U317 ( .A0(R1[6]), .A1(n136), .B0(Rin[6]), .B1(n266), .Y(n421) );
  AOI22X1 U318 ( .A0(L1[2]), .A1(n136), .B0(Lin[2]), .B1(n271), .Y(n479) );
  INVX1 U319 ( .A(n418), .Y(n300) );
  AOI22X1 U320 ( .A0(n194), .A1(n59), .B0(start), .B1(n276), .Y(n418) );
  INVX1 U321 ( .A(n419), .Y(n301) );
  AOI22X1 U322 ( .A0(n63), .A1(n59), .B0(n198), .B1(S2), .Y(n419) );
  INVX1 U323 ( .A(stop_i), .Y(n62) );
endmodule


module euclidean_cell_0 ( deg_Ri, deg_Qi, stop_i, Rin, Qin, Lin, Uin, start, 
        start_cnt, deg_Ro, deg_Qo, stop_o, Rout, Qout, Lout, Uout, st_out, clk, 
        reset );
  input [4:0] deg_Ri;
  input [4:0] deg_Qi;
  input [12:0] Rin;
  input [12:0] Qin;
  input [12:0] Lin;
  input [12:0] Uin;
  output [4:0] deg_Ro;
  output [4:0] deg_Qo;
  output [12:0] Rout;
  output [12:0] Qout;
  output [12:0] Lout;
  output [12:0] Uout;
  input stop_i, start, start_cnt, clk, reset;
  output stop_o, st_out;
  wire   sw, S2, n2, n57, n58, n59, n62, n63, n64, n65, n122, n123, n124, n126,
         n127, n128, n129, n130, n134, n136, n193, n194, n195, n197, n198,
         n199, n200, n201, n258, n259, n260, n262, n263, n264, n265, n266,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535;
  wire   [12:0] d1out;
  wire   [12:0] Q1;
  wire   [12:0] R1;
  wire   [12:0] r_mux;
  wire   [12:0] q_mux;
  wire   [12:0] U1;
  wire   [12:0] L1;
  wire   [12:0] l_mux;
  wire   [12:0] u_mux;
  wire   [12:0] d2out;
  wire   [12:0] d3out;
  wire   [12:0] d4out;
  wire   [12:0] R2;
  wire   [12:0] m1out;
  wire   [12:0] Q2;
  wire   [12:0] m2out;
  wire   [12:0] L2;
  wire   [12:0] m3out;
  wire   [12:0] U2;
  wire   [12:0] m4out;
  wire   [12:0] add1out;
  wire   [12:0] add2out;
  wire   [12:0] Q3;
  wire   [12:0] U3;

  DFFRHQX4 \R2_reg[11]  ( .D(n346), .CK(clk), .RN(reset), .Q(R2[11]) );
  DFFRHQX4 \R2_reg[12]  ( .D(n347), .CK(clk), .RN(reset), .Q(R2[12]) );
  DFFRHQX4 \U2_reg[3]  ( .D(n382), .CK(clk), .RN(reset), .Q(U2[3]) );
  DFFRHQX4 \U2_reg[10]  ( .D(n389), .CK(clk), .RN(reset), .Q(U2[10]) );
  DFFRHQX4 \L2_reg[11]  ( .D(n403), .CK(clk), .RN(reset), .Q(L2[11]) );
  DFFRHQX4 \L2_reg[12]  ( .D(n404), .CK(clk), .RN(reset), .Q(L2[12]) );
  degree_computation_0 degree1 ( .deg_Ri(deg_Ri), .deg_Qi(deg_Qi), .stop_i(n63), .d1out(d1out), .start(start), .deg_Ro(deg_Ro), .deg_Qo(deg_Qo), .stop_o(
        stop_o), .sw(sw), .clk(clk), .reset(reset) );
  mux_13_28 m1 ( .a(Q1), .b(R1), .sel(sw), .out(r_mux) );
  mux_13_27 m2 ( .a(R1), .b(Q1), .sel(sw), .out(q_mux) );
  mux_13_26 m3 ( .a(U1), .b(L1), .sel(sw), .out(l_mux) );
  mux_13_25 m4 ( .a(L1), .b(U1), .sel(sw), .out(u_mux) );
  feedback_ckt_3 D1 ( .Din(q_mux), .start(n2), .Qout(d1out), .clk(clk), 
        .reset(reset) );
  feedback_ckt_2 D2 ( .Din(r_mux), .start(n2), .Qout(d2out), .clk(clk), 
        .reset(reset) );
  feedback_ckt_1 D3 ( .Din(q_mux), .start(n62), .Qout(d3out), .clk(clk), 
        .reset(reset) );
  feedback_ckt_0 D4 ( .Din(r_mux), .start(n62), .Qout(d4out), .clk(clk), 
        .reset(reset) );
  multiplier_3 mx1 ( .a(R2), .b(d1out), .c(m1out) );
  multiplier_2 mx2 ( .a(d2out), .b(Q2), .c(m2out) );
  multiplier_1 mx3 ( .a(L2), .b(d3out), .c(m3out) );
  multiplier_0 mx4 ( .a(d4out), .b(U2), .c(m4out) );
  mux_13_24 m5 ( .a(R2), .b(add1out), .sel(n63), .out(Rout) );
  mux_13_23 m6 ( .a(Q2), .b(Q3), .sel(n63), .out(Qout) );
  mux_13_22 m7 ( .a(L2), .b(add2out), .sel(n63), .out(Lout) );
  mux_13_21 m8 ( .a({U2[12:3], n59, U2[1:0]}), .b(U3), .sel(stop_i), .out(Uout) );
  DFFRHQXL \R1_reg[12]  ( .D(n304), .CK(clk), .RN(reset), .Q(R1[12]) );
  DFFRHQXL \L1_reg[2]  ( .D(n363), .CK(clk), .RN(reset), .Q(L1[2]) );
  DFFSX1 S3_reg ( .D(n418), .CK(clk), .SN(reset), .Q(st_out), .QN(n419) );
  DFFSX1 S2_reg ( .D(n303), .CK(clk), .SN(reset), .Q(S2) );
  DFFRHQX1 \U3_reg[3]  ( .D(n414), .CK(clk), .RN(reset), .Q(U3[3]) );
  DFFRHQX1 \U3_reg[2]  ( .D(n415), .CK(clk), .RN(reset), .Q(U3[2]) );
  DFFRHQX1 \Q3_reg[12]  ( .D(n348), .CK(clk), .RN(reset), .Q(Q3[12]) );
  DFFRHQX1 \Q3_reg[11]  ( .D(n349), .CK(clk), .RN(reset), .Q(Q3[11]) );
  DFFRHQX1 \Q3_reg[10]  ( .D(n350), .CK(clk), .RN(reset), .Q(Q3[10]) );
  DFFRHQX1 \Q3_reg[9]  ( .D(n351), .CK(clk), .RN(reset), .Q(Q3[9]) );
  DFFRHQX1 \Q3_reg[8]  ( .D(n352), .CK(clk), .RN(reset), .Q(Q3[8]) );
  DFFRHQX1 \Q3_reg[7]  ( .D(n353), .CK(clk), .RN(reset), .Q(Q3[7]) );
  DFFRHQX1 \Q3_reg[6]  ( .D(n354), .CK(clk), .RN(reset), .Q(Q3[6]) );
  DFFRHQX1 \Q3_reg[5]  ( .D(n355), .CK(clk), .RN(reset), .Q(Q3[5]) );
  DFFRHQX1 \Q3_reg[4]  ( .D(n356), .CK(clk), .RN(reset), .Q(Q3[4]) );
  DFFRHQX1 \Q3_reg[3]  ( .D(n357), .CK(clk), .RN(reset), .Q(Q3[3]) );
  DFFRHQX1 \Q3_reg[2]  ( .D(n358), .CK(clk), .RN(reset), .Q(Q3[2]) );
  DFFRHQX1 \Q3_reg[1]  ( .D(n359), .CK(clk), .RN(reset), .Q(Q3[1]) );
  DFFRHQX1 \Q3_reg[0]  ( .D(n360), .CK(clk), .RN(reset), .Q(Q3[0]) );
  DFFRHQX1 \U3_reg[12]  ( .D(n405), .CK(clk), .RN(reset), .Q(U3[12]) );
  DFFRHQX1 \U3_reg[11]  ( .D(n406), .CK(clk), .RN(reset), .Q(U3[11]) );
  DFFRHQX1 \U3_reg[10]  ( .D(n407), .CK(clk), .RN(reset), .Q(U3[10]) );
  DFFRHQX1 \U3_reg[9]  ( .D(n408), .CK(clk), .RN(reset), .Q(U3[9]) );
  DFFRHQX1 \U3_reg[8]  ( .D(n409), .CK(clk), .RN(reset), .Q(U3[8]) );
  DFFRHQX1 \U3_reg[7]  ( .D(n410), .CK(clk), .RN(reset), .Q(U3[7]) );
  DFFRHQX1 \U3_reg[6]  ( .D(n411), .CK(clk), .RN(reset), .Q(U3[6]) );
  DFFRHQX1 \U3_reg[5]  ( .D(n412), .CK(clk), .RN(reset), .Q(U3[5]) );
  DFFRHQX1 \U3_reg[4]  ( .D(n413), .CK(clk), .RN(reset), .Q(U3[4]) );
  DFFRHQX1 \U3_reg[1]  ( .D(n416), .CK(clk), .RN(reset), .Q(U3[1]) );
  DFFRHQX1 \U3_reg[0]  ( .D(n417), .CK(clk), .RN(reset), .Q(U3[0]) );
  DFFRHQX1 \R1_reg[1]  ( .D(n307), .CK(clk), .RN(reset), .Q(R1[1]) );
  DFFRHQX1 \R1_reg[0]  ( .D(n308), .CK(clk), .RN(reset), .Q(R1[0]) );
  DFFRHQX1 \Q1_reg[12]  ( .D(n309), .CK(clk), .RN(reset), .Q(Q1[12]) );
  DFFRHQX1 \Q1_reg[11]  ( .D(n310), .CK(clk), .RN(reset), .Q(Q1[11]) );
  DFFRHQX1 \Q1_reg[10]  ( .D(n311), .CK(clk), .RN(reset), .Q(Q1[10]) );
  DFFRHQX1 \Q1_reg[8]  ( .D(n313), .CK(clk), .RN(reset), .Q(Q1[8]) );
  DFFRHQX1 \Q1_reg[7]  ( .D(n314), .CK(clk), .RN(reset), .Q(Q1[7]) );
  DFFRHQX1 \Q1_reg[6]  ( .D(n315), .CK(clk), .RN(reset), .Q(Q1[6]) );
  DFFRHQX1 \Q1_reg[5]  ( .D(n316), .CK(clk), .RN(reset), .Q(Q1[5]) );
  DFFRHQX1 \Q1_reg[4]  ( .D(n317), .CK(clk), .RN(reset), .Q(Q1[4]) );
  DFFRHQX1 \Q1_reg[3]  ( .D(n318), .CK(clk), .RN(reset), .Q(Q1[3]) );
  DFFRHQX1 \Q1_reg[2]  ( .D(n319), .CK(clk), .RN(reset), .Q(Q1[2]) );
  DFFRHQX1 \Q1_reg[1]  ( .D(n320), .CK(clk), .RN(reset), .Q(Q1[1]) );
  DFFRHQX1 \Q1_reg[0]  ( .D(n321), .CK(clk), .RN(reset), .Q(Q1[0]) );
  DFFRHQXL \L1_reg[12]  ( .D(n361), .CK(clk), .RN(reset), .Q(L1[12]) );
  DFFRHQX1 \L1_reg[1]  ( .D(n364), .CK(clk), .RN(reset), .Q(L1[1]) );
  DFFRHQX1 \L1_reg[0]  ( .D(n365), .CK(clk), .RN(reset), .Q(L1[0]) );
  DFFRHQX1 \U1_reg[12]  ( .D(n366), .CK(clk), .RN(reset), .Q(U1[12]) );
  DFFRHQX1 \U1_reg[11]  ( .D(n367), .CK(clk), .RN(reset), .Q(U1[11]) );
  DFFRHQX1 \U1_reg[10]  ( .D(n368), .CK(clk), .RN(reset), .Q(U1[10]) );
  DFFRHQX1 \U1_reg[8]  ( .D(n370), .CK(clk), .RN(reset), .Q(U1[8]) );
  DFFRHQX1 \U1_reg[7]  ( .D(n371), .CK(clk), .RN(reset), .Q(U1[7]) );
  DFFRHQX1 \U1_reg[6]  ( .D(n372), .CK(clk), .RN(reset), .Q(U1[6]) );
  DFFRHQX1 \U1_reg[5]  ( .D(n373), .CK(clk), .RN(reset), .Q(U1[5]) );
  DFFRHQX1 \U1_reg[4]  ( .D(n374), .CK(clk), .RN(reset), .Q(U1[4]) );
  DFFRHQX1 \U1_reg[3]  ( .D(n375), .CK(clk), .RN(reset), .Q(U1[3]) );
  DFFRHQX1 \U1_reg[2]  ( .D(n376), .CK(clk), .RN(reset), .Q(U1[2]) );
  DFFRHQX1 \U1_reg[1]  ( .D(n377), .CK(clk), .RN(reset), .Q(U1[1]) );
  DFFRHQX1 \U1_reg[0]  ( .D(n378), .CK(clk), .RN(reset), .Q(U1[0]) );
  DFFRHQX1 \Q1_reg[9]  ( .D(n312), .CK(clk), .RN(reset), .Q(Q1[9]) );
  DFFRHQX1 \U1_reg[9]  ( .D(n369), .CK(clk), .RN(reset), .Q(U1[9]) );
  DFFRHQX1 \R1_reg[7]  ( .D(n290), .CK(clk), .RN(reset), .Q(R1[7]) );
  DFFRHQX1 \L1_reg[4]  ( .D(n300), .CK(clk), .RN(reset), .Q(L1[4]) );
  DFFRHQX1 \L1_reg[9]  ( .D(n296), .CK(clk), .RN(reset), .Q(L1[9]) );
  DFFSX1 S1_reg ( .D(n302), .CK(clk), .SN(reset), .Q(n2), .QN(n57) );
  DFFRHQX1 \L2_reg[0]  ( .D(n392), .CK(clk), .RN(reset), .Q(L2[0]) );
  DFFRHQX1 \R2_reg[0]  ( .D(n335), .CK(clk), .RN(reset), .Q(R2[0]) );
  DFFRHQX1 \R2_reg[1]  ( .D(n336), .CK(clk), .RN(reset), .Q(R2[1]) );
  DFFRHQX1 \R2_reg[2]  ( .D(n337), .CK(clk), .RN(reset), .Q(R2[2]) );
  DFFRHQX1 \R2_reg[6]  ( .D(n341), .CK(clk), .RN(reset), .Q(R2[6]) );
  DFFRHQX1 \L2_reg[1]  ( .D(n393), .CK(clk), .RN(reset), .Q(L2[1]) );
  DFFRHQX1 \L2_reg[2]  ( .D(n394), .CK(clk), .RN(reset), .Q(L2[2]) );
  DFFRHQX1 \L2_reg[6]  ( .D(n398), .CK(clk), .RN(reset), .Q(L2[6]) );
  DFFRHQX1 \R2_reg[3]  ( .D(n338), .CK(clk), .RN(reset), .Q(R2[3]) );
  DFFRHQX1 \R2_reg[4]  ( .D(n339), .CK(clk), .RN(reset), .Q(R2[4]) );
  DFFRHQX1 \R2_reg[5]  ( .D(n340), .CK(clk), .RN(reset), .Q(R2[5]) );
  DFFRHQX1 \R2_reg[7]  ( .D(n342), .CK(clk), .RN(reset), .Q(R2[7]) );
  DFFRHQX1 \R2_reg[8]  ( .D(n343), .CK(clk), .RN(reset), .Q(R2[8]) );
  DFFRHQX1 \R2_reg[9]  ( .D(n344), .CK(clk), .RN(reset), .Q(R2[9]) );
  DFFRHQX1 \R2_reg[10]  ( .D(n345), .CK(clk), .RN(reset), .Q(R2[10]) );
  DFFRHQX1 \L2_reg[3]  ( .D(n395), .CK(clk), .RN(reset), .Q(L2[3]) );
  DFFRHQX1 \L2_reg[4]  ( .D(n396), .CK(clk), .RN(reset), .Q(L2[4]) );
  DFFRHQX1 \L2_reg[5]  ( .D(n397), .CK(clk), .RN(reset), .Q(L2[5]) );
  DFFRHQX1 \L2_reg[7]  ( .D(n399), .CK(clk), .RN(reset), .Q(L2[7]) );
  DFFRHQX1 \L2_reg[10]  ( .D(n402), .CK(clk), .RN(reset), .Q(L2[10]) );
  DFFRHQX1 \Q2_reg[2]  ( .D(n324), .CK(clk), .RN(reset), .Q(Q2[2]) );
  DFFRHQX1 \Q2_reg[5]  ( .D(n327), .CK(clk), .RN(reset), .Q(Q2[5]) );
  DFFRHQX1 \Q2_reg[6]  ( .D(n328), .CK(clk), .RN(reset), .Q(Q2[6]) );
  DFFRHQX1 \Q2_reg[8]  ( .D(n330), .CK(clk), .RN(reset), .Q(Q2[8]) );
  DFFRHQX1 \Q2_reg[12]  ( .D(n334), .CK(clk), .RN(reset), .Q(Q2[12]) );
  DFFRHQX1 \U2_reg[7]  ( .D(n386), .CK(clk), .RN(reset), .Q(U2[7]) );
  DFFRHQX1 \U2_reg[12]  ( .D(n391), .CK(clk), .RN(reset), .Q(U2[12]) );
  DFFRHQX1 \Q2_reg[9]  ( .D(n331), .CK(clk), .RN(reset), .Q(Q2[9]) );
  DFFRHQX1 \Q2_reg[0]  ( .D(n322), .CK(clk), .RN(reset), .Q(Q2[0]) );
  DFFRHQX1 \U2_reg[0]  ( .D(n379), .CK(clk), .RN(reset), .Q(U2[0]) );
  DFFRHQX1 \Q2_reg[1]  ( .D(n323), .CK(clk), .RN(reset), .Q(Q2[1]) );
  DFFRHQXL \R1_reg[11]  ( .D(n286), .CK(clk), .RN(reset), .Q(R1[11]) );
  DFFRHQXL \R1_reg[10]  ( .D(n287), .CK(clk), .RN(reset), .Q(R1[10]) );
  DFFRHQXL \R1_reg[8]  ( .D(n289), .CK(clk), .RN(reset), .Q(R1[8]) );
  DFFRHQXL \R1_reg[3]  ( .D(n293), .CK(clk), .RN(reset), .Q(R1[3]) );
  DFFRHQXL \L1_reg[11]  ( .D(n294), .CK(clk), .RN(reset), .Q(L1[11]) );
  DFFRHQXL \L1_reg[10]  ( .D(n295), .CK(clk), .RN(reset), .Q(L1[10]) );
  DFFRHQXL \L1_reg[8]  ( .D(n297), .CK(clk), .RN(reset), .Q(L1[8]) );
  DFFRHQXL \L1_reg[7]  ( .D(n298), .CK(clk), .RN(reset), .Q(L1[7]) );
  DFFRHQXL \L1_reg[3]  ( .D(n301), .CK(clk), .RN(reset), .Q(L1[3]) );
  DFFRHQXL \R1_reg[9]  ( .D(n288), .CK(clk), .RN(reset), .Q(R1[9]) );
  DFFRHQXL \R1_reg[4]  ( .D(n292), .CK(clk), .RN(reset), .Q(R1[4]) );
  DFFRHQX4 \U2_reg[2]  ( .D(n381), .CK(clk), .RN(reset), .Q(U2[2]) );
  DFFRHQX1 \U2_reg[5]  ( .D(n384), .CK(clk), .RN(reset), .Q(U2[5]) );
  DFFRHQX2 \Q2_reg[10]  ( .D(n332), .CK(clk), .RN(reset), .Q(Q2[10]) );
  DFFRHQX2 \Q2_reg[11]  ( .D(n333), .CK(clk), .RN(reset), .Q(Q2[11]) );
  DFFRHQXL \L1_reg[5]  ( .D(n299), .CK(clk), .RN(reset), .Q(L1[5]) );
  DFFRHQXL \R1_reg[5]  ( .D(n291), .CK(clk), .RN(reset), .Q(R1[5]) );
  DFFRHQXL \L1_reg[6]  ( .D(n362), .CK(clk), .RN(reset), .Q(L1[6]) );
  DFFRHQXL \R1_reg[6]  ( .D(n305), .CK(clk), .RN(reset), .Q(R1[6]) );
  DFFRHQX2 \Q2_reg[7]  ( .D(n329), .CK(clk), .RN(reset), .Q(Q2[7]) );
  DFFRHQXL \R1_reg[2]  ( .D(n306), .CK(clk), .RN(reset), .Q(R1[2]) );
  DFFRHQX2 \U2_reg[8]  ( .D(n387), .CK(clk), .RN(reset), .Q(U2[8]) );
  DFFRHQX2 \U2_reg[11]  ( .D(n390), .CK(clk), .RN(reset), .Q(U2[11]) );
  DFFRHQX2 \U2_reg[9]  ( .D(n388), .CK(clk), .RN(reset), .Q(U2[9]) );
  DFFRHQX2 \U2_reg[6]  ( .D(n385), .CK(clk), .RN(reset), .Q(U2[6]) );
  DFFRHQX2 \Q2_reg[4]  ( .D(n326), .CK(clk), .RN(reset), .Q(Q2[4]) );
  DFFRHQX2 \Q2_reg[3]  ( .D(n325), .CK(clk), .RN(reset), .Q(Q2[3]) );
  DFFRHQX2 \U2_reg[1]  ( .D(n380), .CK(clk), .RN(reset), .Q(U2[1]) );
  DFFRHQX2 \U2_reg[4]  ( .D(n383), .CK(clk), .RN(reset), .Q(U2[4]) );
  DFFRHQX2 \L2_reg[8]  ( .D(n400), .CK(clk), .RN(reset), .Q(L2[8]) );
  DFFRHQX2 \L2_reg[9]  ( .D(n401), .CK(clk), .RN(reset), .Q(L2[9]) );
  XNOR2X1 U2_inst ( .A(m4out[3]), .B(n279), .Y(add2out[3]) );
  MX2X1 U3_inst ( .A(Rin[5]), .B(R1[5]), .S0(n197), .Y(n291) );
  INVX1 U4 ( .A(L1[12]), .Y(n58) );
  AOI22XL U5 ( .A0(L2[5]), .A1(n199), .B0(l_mux[5]), .B1(n258), .Y(n515) );
  MX2X2 U6 ( .A(Lin[5]), .B(L1[5]), .S0(n195), .Y(n299) );
  AOI2BB2X1 U7 ( .B0(Lin[12]), .B1(n273), .A0N(n58), .A1N(n270), .Y(n479) );
  AOI22X1 U8 ( .A0(Rin[12]), .A1(n271), .B0(R1[12]), .B1(n130), .Y(n422) );
  CLKBUFXL U9 ( .A(U2[2]), .Y(n59) );
  MX2X1 U10 ( .A(R1[7]), .B(Rin[7]), .S0(n258), .Y(n290) );
  XOR2X1 U11 ( .A(m2out[5]), .B(m1out[5]), .Y(add1out[5]) );
  INVXL U12 ( .A(n479), .Y(n361) );
  MX2X1 U13 ( .A(L1[8]), .B(Lin[8]), .S0(n272), .Y(n297) );
  MX2X1 U14 ( .A(L1[7]), .B(Lin[7]), .S0(n274), .Y(n298) );
  MX2X1 U15 ( .A(R1[3]), .B(Rin[3]), .S0(n266), .Y(n293) );
  MX2X1 U16 ( .A(L1[10]), .B(Lin[10]), .S0(n260), .Y(n295) );
  MX2X1 U17 ( .A(L1[3]), .B(Lin[3]), .S0(n270), .Y(n301) );
  MX2X1 U18 ( .A(L1[4]), .B(Lin[4]), .S0(n275), .Y(n300) );
  MX2X1 U19 ( .A(L1[11]), .B(Lin[11]), .S0(n274), .Y(n294) );
  MX2X1 U20 ( .A(R1[8]), .B(Rin[8]), .S0(n275), .Y(n289) );
  MX2X1 U21 ( .A(R1[10]), .B(Rin[10]), .S0(n270), .Y(n287) );
  MX2X1 U22 ( .A(R1[11]), .B(Rin[11]), .S0(n274), .Y(n286) );
  MX2X1 U23 ( .A(R1[9]), .B(Rin[9]), .S0(n266), .Y(n288) );
  INVXL U24 ( .A(n422), .Y(n304) );
  INVXL U25 ( .A(n481), .Y(n363) );
  INVXL U26 ( .A(n423), .Y(n305) );
  INVXL U27 ( .A(n425), .Y(n307) );
  INVXL U28 ( .A(n424), .Y(n306) );
  INVXL U29 ( .A(n482), .Y(n364) );
  INVXL U30 ( .A(n480), .Y(n362) );
  AOI22XL U31 ( .A0(n266), .A1(n59), .B0(U3[2]), .B1(n200), .Y(n533) );
  AOI22XL U32 ( .A0(n258), .A1(Q2[1]), .B0(Q3[1]), .B1(n199), .Y(n477) );
  AOI22XL U33 ( .A0(L2[12]), .A1(n129), .B0(l_mux[12]), .B1(n273), .Y(n522) );
  AOI22XL U34 ( .A0(L2[11]), .A1(n194), .B0(l_mux[11]), .B1(n270), .Y(n521) );
  AOI22XL U35 ( .A0(n198), .A1(U2[11]), .B0(u_mux[11]), .B1(n65), .Y(n508) );
  AOI22XL U36 ( .A0(n277), .A1(U2[10]), .B0(u_mux[10]), .B1(n264), .Y(n507) );
  AOI22XL U37 ( .A0(n197), .A1(U2[9]), .B0(u_mux[9]), .B1(n260), .Y(n506) );
  AOI22XL U38 ( .A0(n195), .A1(U2[6]), .B0(u_mux[6]), .B1(n260), .Y(n503) );
  AOI22XL U39 ( .A0(n193), .A1(U2[4]), .B0(u_mux[4]), .B1(n259), .Y(n501) );
  AOI22XL U40 ( .A0(n194), .A1(U2[3]), .B0(u_mux[3]), .B1(n264), .Y(n500) );
  AOI22XL U41 ( .A0(n128), .A1(U2[1]), .B0(u_mux[1]), .B1(n266), .Y(n498) );
  AOI22XL U42 ( .A0(R2[12]), .A1(n197), .B0(r_mux[12]), .B1(n264), .Y(n465) );
  AOI22XL U43 ( .A0(R2[11]), .A1(n127), .B0(r_mux[11]), .B1(n274), .Y(n464) );
  AOI22XL U44 ( .A0(n136), .A1(Q2[11]), .B0(q_mux[11]), .B1(n65), .Y(n451) );
  AOI22XL U45 ( .A0(n128), .A1(Q2[3]), .B0(q_mux[3]), .B1(n258), .Y(n443) );
  AOI22XL U46 ( .A0(n271), .A1(U2[0]), .B0(U3[0]), .B1(n199), .Y(n535) );
  AOI22XL U47 ( .A0(n273), .A1(U2[1]), .B0(U3[1]), .B1(n278), .Y(n534) );
  AOI22XL U48 ( .A0(n194), .A1(n59), .B0(u_mux[2]), .B1(n265), .Y(n499) );
  AOI22XL U49 ( .A0(L2[9]), .A1(n199), .B0(l_mux[9]), .B1(n274), .Y(n519) );
  AOI22XL U50 ( .A0(L2[8]), .A1(n194), .B0(l_mux[8]), .B1(n258), .Y(n518) );
  AOI22XL U51 ( .A0(L2[3]), .A1(n136), .B0(l_mux[3]), .B1(n272), .Y(n513) );
  AOI22XL U52 ( .A0(n278), .A1(U2[12]), .B0(u_mux[12]), .B1(n265), .Y(n509) );
  AOI22XL U53 ( .A0(n130), .A1(U2[8]), .B0(u_mux[8]), .B1(n273), .Y(n505) );
  AOI22XL U54 ( .A0(n197), .A1(U2[7]), .B0(u_mux[7]), .B1(n262), .Y(n504) );
  AOI22XL U55 ( .A0(n195), .A1(U2[5]), .B0(u_mux[5]), .B1(n272), .Y(n502) );
  AOI22XL U56 ( .A0(n195), .A1(U2[0]), .B0(u_mux[0]), .B1(n273), .Y(n497) );
  AOI22XL U57 ( .A0(R2[10]), .A1(n128), .B0(r_mux[10]), .B1(n274), .Y(n463) );
  AOI22XL U58 ( .A0(R2[9]), .A1(n127), .B0(r_mux[9]), .B1(n259), .Y(n462) );
  AOI22XL U59 ( .A0(R2[8]), .A1(n194), .B0(r_mux[8]), .B1(n260), .Y(n461) );
  AOI22XL U60 ( .A0(R2[7]), .A1(n200), .B0(r_mux[7]), .B1(n258), .Y(n460) );
  AOI22XL U61 ( .A0(R2[6]), .A1(n278), .B0(r_mux[6]), .B1(n263), .Y(n459) );
  AOI22XL U62 ( .A0(R2[5]), .A1(n201), .B0(r_mux[5]), .B1(n274), .Y(n458) );
  AOI22XL U63 ( .A0(R2[4]), .A1(n198), .B0(r_mux[4]), .B1(n275), .Y(n457) );
  AOI22XL U64 ( .A0(R2[3]), .A1(n199), .B0(r_mux[3]), .B1(n65), .Y(n456) );
  AOI22XL U65 ( .A0(n130), .A1(Q2[12]), .B0(q_mux[12]), .B1(n271), .Y(n452) );
  AOI22XL U66 ( .A0(n136), .A1(Q2[9]), .B0(q_mux[9]), .B1(n271), .Y(n449) );
  AOI22XL U67 ( .A0(n194), .A1(Q2[8]), .B0(q_mux[8]), .B1(n265), .Y(n448) );
  AOI22XL U68 ( .A0(n129), .A1(Q2[7]), .B0(q_mux[7]), .B1(n259), .Y(n447) );
  AOI22XL U69 ( .A0(n134), .A1(Q2[6]), .B0(q_mux[6]), .B1(n273), .Y(n446) );
  AOI22XL U70 ( .A0(n129), .A1(Q2[5]), .B0(q_mux[5]), .B1(n259), .Y(n445) );
  AOI22XL U71 ( .A0(n134), .A1(Q2[4]), .B0(q_mux[4]), .B1(n260), .Y(n444) );
  AOI22XL U72 ( .A0(n128), .A1(Q2[1]), .B0(q_mux[1]), .B1(n259), .Y(n441) );
  AOI22XL U73 ( .A0(n130), .A1(Q2[0]), .B0(q_mux[0]), .B1(n258), .Y(n440) );
  AOI22XL U74 ( .A0(n122), .A1(U2[3]), .B0(U3[3]), .B1(n276), .Y(n532) );
  AOI22XL U75 ( .A0(n274), .A1(U2[4]), .B0(U3[4]), .B1(n200), .Y(n531) );
  AOI22XL U76 ( .A0(n275), .A1(U2[5]), .B0(U3[5]), .B1(n201), .Y(n530) );
  AOI22XL U77 ( .A0(n270), .A1(U2[6]), .B0(U3[6]), .B1(n199), .Y(n529) );
  AOI22XL U78 ( .A0(n266), .A1(U2[7]), .B0(U3[7]), .B1(n201), .Y(n528) );
  AOI22XL U79 ( .A0(n274), .A1(U2[8]), .B0(U3[8]), .B1(n201), .Y(n527) );
  AOI22XL U80 ( .A0(n271), .A1(U2[9]), .B0(U3[9]), .B1(n201), .Y(n526) );
  AOI22XL U81 ( .A0(n122), .A1(U2[10]), .B0(U3[10]), .B1(n277), .Y(n525) );
  AOI22XL U82 ( .A0(n272), .A1(U2[11]), .B0(U3[11]), .B1(n201), .Y(n524) );
  AOI22XL U83 ( .A0(n271), .A1(U2[12]), .B0(U3[12]), .B1(n201), .Y(n523) );
  AOI22XL U84 ( .A0(n270), .A1(Q2[0]), .B0(Q3[0]), .B1(n199), .Y(n478) );
  AOI22XL U85 ( .A0(n273), .A1(Q2[3]), .B0(Q3[3]), .B1(n277), .Y(n475) );
  AOI22XL U86 ( .A0(n272), .A1(Q2[4]), .B0(Q3[4]), .B1(n276), .Y(n474) );
  AOI22XL U87 ( .A0(n275), .A1(Q2[5]), .B0(Q3[5]), .B1(n198), .Y(n473) );
  AOI22XL U88 ( .A0(n258), .A1(Q2[6]), .B0(Q3[6]), .B1(n200), .Y(n472) );
  AOI22XL U89 ( .A0(n271), .A1(Q2[9]), .B0(Q3[9]), .B1(n276), .Y(n469) );
  AOI22XL U90 ( .A0(n266), .A1(Q2[12]), .B0(Q3[12]), .B1(n201), .Y(n466) );
  AOI22XL U91 ( .A0(n266), .A1(Q2[7]), .B0(Q3[7]), .B1(n276), .Y(n471) );
  AOI22XL U92 ( .A0(n275), .A1(Q2[8]), .B0(Q3[8]), .B1(n200), .Y(n470) );
  AOI22XL U93 ( .A0(n273), .A1(Q2[11]), .B0(Q3[11]), .B1(n278), .Y(n467) );
  INVX1 U94 ( .A(n265), .Y(n124) );
  INVX1 U95 ( .A(n265), .Y(n126) );
  INVX1 U96 ( .A(n264), .Y(n127) );
  INVX1 U97 ( .A(n260), .Y(n197) );
  INVX1 U98 ( .A(n260), .Y(n195) );
  INVX1 U99 ( .A(n266), .Y(n194) );
  INVX1 U100 ( .A(n262), .Y(n193) );
  INVX1 U101 ( .A(n263), .Y(n136) );
  INVX1 U102 ( .A(n264), .Y(n129) );
  INVX1 U103 ( .A(n263), .Y(n134) );
  INVX1 U104 ( .A(n264), .Y(n128) );
  INVX1 U105 ( .A(n263), .Y(n130) );
  INVX1 U106 ( .A(n260), .Y(n198) );
  INVX1 U107 ( .A(n259), .Y(n201) );
  INVX1 U108 ( .A(n65), .Y(n199) );
  INVX1 U109 ( .A(n65), .Y(n200) );
  INVX1 U110 ( .A(n278), .Y(n259) );
  INVX1 U111 ( .A(n276), .Y(n265) );
  INVX1 U112 ( .A(n277), .Y(n260) );
  INVX1 U113 ( .A(n123), .Y(n272) );
  INVX1 U114 ( .A(n123), .Y(n266) );
  INVX1 U115 ( .A(n276), .Y(n271) );
  INVX1 U116 ( .A(n278), .Y(n270) );
  INVX1 U117 ( .A(n123), .Y(n273) );
  INVX1 U118 ( .A(n277), .Y(n262) );
  INVX1 U119 ( .A(n276), .Y(n264) );
  INVX1 U120 ( .A(n276), .Y(n263) );
  INVX1 U121 ( .A(n123), .Y(n274) );
  INVX1 U122 ( .A(n277), .Y(n275) );
  INVX1 U123 ( .A(n123), .Y(n258) );
  INVX1 U124 ( .A(n122), .Y(n278) );
  INVX1 U125 ( .A(n122), .Y(n276) );
  INVX1 U126 ( .A(n122), .Y(n277) );
  INVX1 U127 ( .A(n123), .Y(n65) );
  INVX1 U128 ( .A(n123), .Y(n122) );
  INVX1 U129 ( .A(start_cnt), .Y(n123) );
  XOR2X1 U130 ( .A(m1out[8]), .B(m2out[8]), .Y(add1out[8]) );
  XOR2X1 U131 ( .A(m1out[4]), .B(m2out[4]), .Y(add1out[4]) );
  XOR2X1 U132 ( .A(m1out[3]), .B(m2out[3]), .Y(add1out[3]) );
  XOR2X1 U133 ( .A(m1out[11]), .B(m2out[11]), .Y(add1out[11]) );
  XOR2X1 U134 ( .A(m1out[10]), .B(m2out[10]), .Y(add1out[10]) );
  XOR2X1 U135 ( .A(m1out[9]), .B(m2out[9]), .Y(add1out[9]) );
  XOR2X1 U136 ( .A(m1out[7]), .B(m2out[7]), .Y(add1out[7]) );
  XOR2X1 U137 ( .A(m2out[6]), .B(m1out[6]), .Y(add1out[6]) );
  XOR2X1 U138 ( .A(m2out[2]), .B(m1out[2]), .Y(add1out[2]) );
  XOR2X1 U139 ( .A(m2out[1]), .B(m1out[1]), .Y(add1out[1]) );
  XOR2X1 U140 ( .A(m2out[12]), .B(m1out[12]), .Y(add1out[12]) );
  INVX1 U141 ( .A(m3out[5]), .Y(n280) );
  INVX1 U142 ( .A(m3out[8]), .Y(n281) );
  INVX1 U143 ( .A(m3out[3]), .Y(n279) );
  XOR2X1 U144 ( .A(m2out[0]), .B(m1out[0]), .Y(add1out[0]) );
  INVX1 U145 ( .A(n57), .Y(n62) );
  INVX1 U146 ( .A(n64), .Y(n63) );
  XNOR2X1 U147 ( .A(m4out[8]), .B(n281), .Y(add2out[8]) );
  XOR2X1 U148 ( .A(m3out[7]), .B(m4out[7]), .Y(add2out[7]) );
  XNOR2X1 U149 ( .A(m4out[5]), .B(n280), .Y(add2out[5]) );
  XOR2X1 U150 ( .A(m3out[10]), .B(m4out[10]), .Y(add2out[10]) );
  XOR2X1 U151 ( .A(m3out[9]), .B(m4out[9]), .Y(add2out[9]) );
  XOR2X1 U152 ( .A(m3out[11]), .B(m4out[11]), .Y(add2out[11]) );
  XOR2X1 U153 ( .A(m3out[4]), .B(m4out[4]), .Y(add2out[4]) );
  MXI2X1 U154 ( .A(n283), .B(n282), .S0(n272), .Y(n296) );
  INVX1 U155 ( .A(L1[9]), .Y(n283) );
  INVX1 U156 ( .A(Lin[9]), .Y(n282) );
  MXI2X1 U157 ( .A(n285), .B(n284), .S0(n263), .Y(n292) );
  INVX1 U158 ( .A(R1[4]), .Y(n285) );
  INVX1 U159 ( .A(Rin[4]), .Y(n284) );
  OAI2BB2X1 U160 ( .B0(n271), .B1(n419), .A0N(S2), .A1N(n272), .Y(n418) );
  XOR2X1 U161 ( .A(m4out[12]), .B(m3out[12]), .Y(add2out[12]) );
  XOR2X1 U162 ( .A(m4out[6]), .B(m3out[6]), .Y(add2out[6]) );
  XOR2X1 U163 ( .A(m4out[2]), .B(m3out[2]), .Y(add2out[2]) );
  XOR2X1 U164 ( .A(m4out[1]), .B(m3out[1]), .Y(add2out[1]) );
  XOR2X1 U165 ( .A(m4out[0]), .B(m3out[0]), .Y(add2out[0]) );
  INVX1 U166 ( .A(n533), .Y(n415) );
  INVX1 U167 ( .A(n532), .Y(n414) );
  AOI22X1 U168 ( .A0(L1[2]), .A1(n126), .B0(Lin[2]), .B1(n260), .Y(n481) );
  INVX1 U169 ( .A(n477), .Y(n359) );
  INVX1 U170 ( .A(n441), .Y(n323) );
  INVX1 U171 ( .A(n534), .Y(n416) );
  INVX1 U172 ( .A(n498), .Y(n380) );
  INVX1 U173 ( .A(n535), .Y(n417) );
  INVX1 U174 ( .A(n497), .Y(n379) );
  INVX1 U175 ( .A(n478), .Y(n360) );
  INVX1 U176 ( .A(n440), .Y(n322) );
  INVX1 U177 ( .A(n526), .Y(n408) );
  INVX1 U178 ( .A(n506), .Y(n388) );
  INVX1 U179 ( .A(n469), .Y(n351) );
  INVX1 U180 ( .A(n449), .Y(n331) );
  INVX1 U181 ( .A(n531), .Y(n413) );
  INVX1 U182 ( .A(n530), .Y(n412) );
  INVX1 U183 ( .A(n529), .Y(n411) );
  INVX1 U184 ( .A(n528), .Y(n410) );
  INVX1 U185 ( .A(n527), .Y(n409) );
  INVX1 U186 ( .A(n525), .Y(n407) );
  INVX1 U187 ( .A(n524), .Y(n406) );
  INVX1 U188 ( .A(n523), .Y(n405) );
  INVX1 U189 ( .A(n509), .Y(n391) );
  INVX1 U190 ( .A(n508), .Y(n390) );
  INVX1 U191 ( .A(n507), .Y(n389) );
  INVX1 U192 ( .A(n505), .Y(n387) );
  INVX1 U193 ( .A(n504), .Y(n386) );
  INVX1 U194 ( .A(n503), .Y(n385) );
  INVX1 U195 ( .A(n502), .Y(n384) );
  INVX1 U196 ( .A(n501), .Y(n383) );
  INVX1 U197 ( .A(n476), .Y(n358) );
  AOI22X1 U198 ( .A0(n258), .A1(Q2[2]), .B0(Q3[2]), .B1(n277), .Y(n476) );
  INVX1 U199 ( .A(n475), .Y(n357) );
  INVX1 U200 ( .A(n474), .Y(n356) );
  INVX1 U201 ( .A(n473), .Y(n355) );
  INVX1 U202 ( .A(n472), .Y(n354) );
  INVX1 U203 ( .A(n471), .Y(n353) );
  INVX1 U204 ( .A(n470), .Y(n352) );
  INVX1 U205 ( .A(n468), .Y(n350) );
  AOI22X1 U206 ( .A0(n122), .A1(Q2[10]), .B0(Q3[10]), .B1(n200), .Y(n468) );
  INVX1 U207 ( .A(n467), .Y(n349) );
  INVX1 U208 ( .A(n466), .Y(n348) );
  INVX1 U209 ( .A(n452), .Y(n334) );
  INVX1 U210 ( .A(n451), .Y(n333) );
  INVX1 U211 ( .A(n450), .Y(n332) );
  AOI22X1 U212 ( .A0(n193), .A1(Q2[10]), .B0(q_mux[10]), .B1(n263), .Y(n450)
         );
  INVX1 U213 ( .A(n448), .Y(n330) );
  INVX1 U214 ( .A(n447), .Y(n329) );
  INVX1 U215 ( .A(n446), .Y(n328) );
  INVX1 U216 ( .A(n445), .Y(n327) );
  INVX1 U217 ( .A(n444), .Y(n326) );
  INVX1 U218 ( .A(n443), .Y(n325) );
  INVX1 U219 ( .A(n442), .Y(n324) );
  AOI22X1 U220 ( .A0(n193), .A1(Q2[2]), .B0(q_mux[2]), .B1(n262), .Y(n442) );
  INVX1 U221 ( .A(n499), .Y(n381) );
  INVX1 U222 ( .A(n519), .Y(n401) );
  INVX1 U223 ( .A(n518), .Y(n400) );
  INVX1 U224 ( .A(n517), .Y(n399) );
  AOI22X1 U225 ( .A0(L2[7]), .A1(n195), .B0(l_mux[7]), .B1(n65), .Y(n517) );
  INVX1 U226 ( .A(n516), .Y(n398) );
  AOI22X1 U227 ( .A0(L2[6]), .A1(n197), .B0(l_mux[6]), .B1(n259), .Y(n516) );
  INVX1 U228 ( .A(n515), .Y(n397) );
  INVX1 U229 ( .A(n514), .Y(n396) );
  AOI22X1 U230 ( .A0(L2[4]), .A1(n193), .B0(l_mux[4]), .B1(n260), .Y(n514) );
  INVX1 U231 ( .A(n513), .Y(n395) );
  INVX1 U232 ( .A(n512), .Y(n394) );
  AOI22X1 U233 ( .A0(L2[2]), .A1(n193), .B0(l_mux[2]), .B1(n262), .Y(n512) );
  INVX1 U234 ( .A(n511), .Y(n393) );
  AOI22X1 U235 ( .A0(L2[1]), .A1(n128), .B0(l_mux[1]), .B1(n270), .Y(n511) );
  INVX1 U236 ( .A(n510), .Y(n392) );
  AOI22X1 U237 ( .A0(L2[0]), .A1(n276), .B0(l_mux[0]), .B1(n262), .Y(n510) );
  INVX1 U238 ( .A(n500), .Y(n382) );
  INVX1 U239 ( .A(n496), .Y(n378) );
  AOI22X1 U240 ( .A0(U1[0]), .A1(n127), .B0(Uin[0]), .B1(n262), .Y(n496) );
  INVX1 U241 ( .A(n495), .Y(n377) );
  AOI22X1 U242 ( .A0(U1[1]), .A1(n193), .B0(Uin[1]), .B1(n263), .Y(n495) );
  INVX1 U243 ( .A(n494), .Y(n376) );
  AOI22X1 U244 ( .A0(U1[2]), .A1(n136), .B0(Uin[2]), .B1(n259), .Y(n494) );
  INVX1 U245 ( .A(n493), .Y(n375) );
  AOI22X1 U246 ( .A0(U1[3]), .A1(n194), .B0(Uin[3]), .B1(n265), .Y(n493) );
  INVX1 U247 ( .A(n492), .Y(n374) );
  AOI22X1 U248 ( .A0(U1[4]), .A1(n129), .B0(Uin[4]), .B1(n264), .Y(n492) );
  INVX1 U249 ( .A(n491), .Y(n373) );
  AOI22X1 U250 ( .A0(U1[5]), .A1(n124), .B0(Uin[5]), .B1(n272), .Y(n491) );
  INVX1 U251 ( .A(n490), .Y(n372) );
  AOI22X1 U252 ( .A0(U1[6]), .A1(n124), .B0(Uin[6]), .B1(n263), .Y(n490) );
  INVX1 U253 ( .A(n489), .Y(n371) );
  AOI22X1 U254 ( .A0(U1[7]), .A1(n127), .B0(Uin[7]), .B1(n65), .Y(n489) );
  INVX1 U255 ( .A(n488), .Y(n370) );
  AOI22X1 U256 ( .A0(U1[8]), .A1(n124), .B0(Uin[8]), .B1(n264), .Y(n488) );
  INVX1 U257 ( .A(n487), .Y(n369) );
  AOI22X1 U258 ( .A0(U1[9]), .A1(n124), .B0(Uin[9]), .B1(n262), .Y(n487) );
  INVX1 U259 ( .A(n486), .Y(n368) );
  AOI22X1 U260 ( .A0(U1[10]), .A1(n124), .B0(Uin[10]), .B1(n263), .Y(n486) );
  INVX1 U261 ( .A(n485), .Y(n367) );
  AOI22X1 U262 ( .A0(U1[11]), .A1(n199), .B0(Uin[11]), .B1(n265), .Y(n485) );
  INVX1 U263 ( .A(n484), .Y(n366) );
  AOI22X1 U264 ( .A0(U1[12]), .A1(n124), .B0(Uin[12]), .B1(n65), .Y(n484) );
  INVX1 U265 ( .A(n483), .Y(n365) );
  AOI22X1 U266 ( .A0(L1[0]), .A1(n126), .B0(Lin[0]), .B1(n65), .Y(n483) );
  AOI22X1 U267 ( .A0(L1[1]), .A1(n126), .B0(Lin[1]), .B1(n65), .Y(n482) );
  INVX1 U268 ( .A(n465), .Y(n347) );
  INVX1 U269 ( .A(n464), .Y(n346) );
  INVX1 U270 ( .A(n463), .Y(n345) );
  INVX1 U271 ( .A(n462), .Y(n344) );
  INVX1 U272 ( .A(n461), .Y(n343) );
  INVX1 U273 ( .A(n460), .Y(n342) );
  INVX1 U274 ( .A(n459), .Y(n341) );
  INVX1 U275 ( .A(n458), .Y(n340) );
  INVX1 U276 ( .A(n457), .Y(n339) );
  INVX1 U277 ( .A(n456), .Y(n338) );
  INVX1 U278 ( .A(n455), .Y(n337) );
  AOI22X1 U279 ( .A0(R2[2]), .A1(n200), .B0(r_mux[2]), .B1(n264), .Y(n455) );
  INVX1 U280 ( .A(n454), .Y(n336) );
  AOI22X1 U281 ( .A0(R2[1]), .A1(n200), .B0(r_mux[1]), .B1(n265), .Y(n454) );
  INVX1 U282 ( .A(n453), .Y(n335) );
  AOI22X1 U283 ( .A0(R2[0]), .A1(n199), .B0(r_mux[0]), .B1(n264), .Y(n453) );
  INVX1 U284 ( .A(n439), .Y(n321) );
  AOI22X1 U285 ( .A0(Q1[0]), .A1(n198), .B0(Qin[0]), .B1(n270), .Y(n439) );
  INVX1 U286 ( .A(n438), .Y(n320) );
  AOI22X1 U287 ( .A0(Q1[1]), .A1(n194), .B0(Qin[1]), .B1(n271), .Y(n438) );
  INVX1 U288 ( .A(n437), .Y(n319) );
  AOI22X1 U289 ( .A0(Q1[2]), .A1(n200), .B0(Qin[2]), .B1(n275), .Y(n437) );
  INVX1 U290 ( .A(n436), .Y(n318) );
  AOI22X1 U291 ( .A0(Q1[3]), .A1(n201), .B0(Qin[3]), .B1(n265), .Y(n436) );
  INVX1 U292 ( .A(n435), .Y(n317) );
  AOI22X1 U293 ( .A0(Q1[4]), .A1(n199), .B0(Qin[4]), .B1(n273), .Y(n435) );
  INVX1 U294 ( .A(n434), .Y(n316) );
  AOI22X1 U295 ( .A0(Q1[5]), .A1(n127), .B0(Qin[5]), .B1(n258), .Y(n434) );
  INVX1 U296 ( .A(n433), .Y(n315) );
  AOI22X1 U297 ( .A0(Q1[6]), .A1(n201), .B0(Qin[6]), .B1(n262), .Y(n433) );
  INVX1 U298 ( .A(n432), .Y(n314) );
  AOI22X1 U299 ( .A0(Q1[7]), .A1(n195), .B0(Qin[7]), .B1(n266), .Y(n432) );
  INVX1 U300 ( .A(n431), .Y(n313) );
  AOI22X1 U301 ( .A0(Q1[8]), .A1(n197), .B0(Qin[8]), .B1(n275), .Y(n431) );
  INVX1 U302 ( .A(n430), .Y(n312) );
  AOI22X1 U303 ( .A0(Q1[9]), .A1(n126), .B0(Qin[9]), .B1(n272), .Y(n430) );
  INVX1 U304 ( .A(n429), .Y(n311) );
  AOI22X1 U305 ( .A0(Q1[10]), .A1(n193), .B0(Qin[10]), .B1(n270), .Y(n429) );
  INVX1 U306 ( .A(n428), .Y(n310) );
  AOI22X1 U307 ( .A0(Q1[11]), .A1(n134), .B0(Qin[11]), .B1(n122), .Y(n428) );
  INVX1 U308 ( .A(n427), .Y(n309) );
  AOI22X1 U309 ( .A0(Q1[12]), .A1(n126), .B0(Qin[12]), .B1(n263), .Y(n427) );
  INVX1 U310 ( .A(n426), .Y(n308) );
  AOI22X1 U311 ( .A0(R1[0]), .A1(n193), .B0(Rin[0]), .B1(n270), .Y(n426) );
  AOI22X1 U312 ( .A0(R1[1]), .A1(n200), .B0(Rin[1]), .B1(n272), .Y(n425) );
  AOI22X1 U313 ( .A0(R1[6]), .A1(n194), .B0(Rin[6]), .B1(n274), .Y(n423) );
  AOI22X1 U314 ( .A0(L1[6]), .A1(n126), .B0(Lin[6]), .B1(n275), .Y(n480) );
  INVX1 U315 ( .A(n522), .Y(n404) );
  INVX1 U316 ( .A(n521), .Y(n403) );
  INVX1 U317 ( .A(n520), .Y(n402) );
  AOI22X1 U318 ( .A0(L2[10]), .A1(n194), .B0(l_mux[10]), .B1(n266), .Y(n520)
         );
  INVX1 U319 ( .A(stop_i), .Y(n64) );
  AOI22X1 U320 ( .A0(R1[2]), .A1(n129), .B0(Rin[2]), .B1(n271), .Y(n424) );
  INVX1 U321 ( .A(n420), .Y(n302) );
  AOI22X1 U322 ( .A0(n134), .A1(n62), .B0(start), .B1(n275), .Y(n420) );
  INVX1 U323 ( .A(n421), .Y(n303) );
  AOI22X1 U324 ( .A0(n273), .A1(n62), .B0(n129), .B1(S2), .Y(n421) );
endmodule


module mux_5_23 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n8, n9, n10, n11, n12, n13;

  INVX1 U1 ( .A(sel), .Y(n9) );
  INVX1 U2 ( .A(n13), .Y(out[0]) );
  AOI22X1 U3 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n9), .Y(n13) );
  INVX1 U4 ( .A(n12), .Y(out[1]) );
  AOI22X1 U5 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n9), .Y(n12) );
  INVX1 U6 ( .A(n11), .Y(out[2]) );
  AOI22X1 U7 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n9), .Y(n11) );
  INVX1 U8 ( .A(n10), .Y(out[3]) );
  AOI22X1 U9 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n9), .Y(n10) );
  INVX1 U10 ( .A(n8), .Y(out[4]) );
  AOI22X1 U11 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n9), .Y(n8) );
endmodule


module multiplier_15 ( a, b, c );
  input [12:0] a;
  input [12:0] b;
  output [12:0] c;
  wire   n40, n41, n42, n43, n44, n45, n46, n48, n56, n69, n70, n71, n72, n73,
         n74, n75, n76, n88, n89, n90, n91, n93, n94, n112, n113, n114, n115,
         n116, n117, n118, n120, n121, n123, n124, n125, n156, n157, n158,
         n159, n160, n161, n171, n172, n183, n184, n185, n186, n197, n198,
         n199, n200, n201, n206, n207, n208, n209, n218, n229, n231, n232,
         n241, n242, n243, n244, n245, n255, n256, n257, n258, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n279, n280,
         n281, n282, n283, n284, n285, n287, n292, n293, n294, n295, n307,
         n308, n309, n310, n312, n313, n328, n340, n341, n342, n344, n345,
         n379, n390, n391, n392, n393, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n47, n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n92, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n119, n122,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n202, n203, n204, n205, n210, n211, n212,
         n213, n214, n215, n216, n217, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n230, n233, n234, n235, n236, n237, n238,
         n239, n240, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n259, n260, n261, n262, n263, n264, n265, n266, n278, n286, n288,
         n289, n290, n291, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n311, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n343, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n394, n395;

  NAND3X1 U1 ( .A(n327), .B(n326), .C(n325), .Y(n386) );
  OAI21XL U2 ( .A0(n382), .A1(n145), .B0(n95), .Y(n146) );
  OAI21XL U3 ( .A0(n1), .A1(n100), .B0(n381), .Y(n252) );
  INVX1 U4 ( .A(n50), .Y(n1) );
  OAI211X1 U5 ( .A0(n378), .A1(n62), .B0(n384), .C0(n383), .Y(n385) );
  OAI21XL U6 ( .A0(n2), .A1(n101), .B0(n317), .Y(n319) );
  INVX1 U7 ( .A(n49), .Y(n2) );
  OAI21XL U8 ( .A0(n382), .A1(n108), .B0(n101), .Y(n109) );
  INVX1 U9 ( .A(n317), .Y(n382) );
  XOR2X2 U10 ( .A(n119), .B(n111), .Y(n376) );
  XOR2X1 U11 ( .A(n386), .B(n6), .Y(n363) );
  NOR2X1 U12 ( .A(n190), .B(n191), .Y(n3) );
  INVX1 U13 ( .A(n3), .Y(n192) );
  NOR2X1 U14 ( .A(n73), .B(n20), .Y(n198) );
  OR2X2 U15 ( .A(n191), .B(n187), .Y(n194) );
  OAI21XL U16 ( .A0(n4), .A1(n323), .B0(n324), .Y(n325) );
  INVX1 U17 ( .A(n322), .Y(n4) );
  NAND3X1 U18 ( .A(n191), .B(n187), .C(n190), .Y(n193) );
  AND2X2 U19 ( .A(n95), .B(n105), .Y(n118) );
  AOI211X1 U20 ( .A0(n319), .A1(n38), .B0(n324), .C0(n39), .Y(n5) );
  INVX1 U21 ( .A(n5), .Y(n327) );
  XNOR2X1 U22 ( .A(n223), .B(n245), .Y(c[1]) );
  XOR2X2 U23 ( .A(n264), .B(n68), .Y(n286) );
  NAND2BX1 U24 ( .AN(a[11]), .B(a[12]), .Y(n317) );
  XOR2X1 U25 ( .A(n162), .B(n155), .Y(n177) );
  NAND2X1 U26 ( .A(n107), .B(n18), .Y(n258) );
  XOR2X4 U27 ( .A(n265), .B(n176), .Y(n204) );
  AOI22XL U28 ( .A0(a[4]), .A1(n160), .B0(a[5]), .B1(n161), .Y(n159) );
  OAI2BB1X1 U29 ( .A0N(a[11]), .A1N(n321), .B0(n92), .Y(n110) );
  XOR2X1 U30 ( .A(n204), .B(n177), .Y(n79) );
  XNOR3X2 U31 ( .A(n54), .B(n55), .C(n302), .Y(n6) );
  AND2X2 U32 ( .A(n104), .B(n38), .Y(n7) );
  XNOR3X2 U33 ( .A(n240), .B(n239), .C(n238), .Y(n8) );
  INVX1 U34 ( .A(n324), .Y(n320) );
  NAND2X1 U35 ( .A(b[1]), .B(n46), .Y(n9) );
  INVX1 U36 ( .A(n216), .Y(n10) );
  INVX1 U37 ( .A(n389), .Y(n11) );
  INVX1 U38 ( .A(b[12]), .Y(n12) );
  INVX1 U39 ( .A(n12), .Y(n13) );
  INVX1 U40 ( .A(n12), .Y(n14) );
  INVX1 U41 ( .A(n166), .Y(n15) );
  INVX1 U42 ( .A(n227), .Y(n16) );
  INVX1 U43 ( .A(b[8]), .Y(n17) );
  INVX1 U44 ( .A(n17), .Y(n18) );
  INVX1 U45 ( .A(n122), .Y(n19) );
  INVX1 U46 ( .A(a[1]), .Y(n20) );
  INVX1 U47 ( .A(n20), .Y(n21) );
  INVX1 U48 ( .A(n56), .Y(n22) );
  INVX1 U49 ( .A(a[3]), .Y(n23) );
  INVXL U50 ( .A(n23), .Y(n24) );
  INVX1 U51 ( .A(a[7]), .Y(n25) );
  INVXL U52 ( .A(n25), .Y(n26) );
  INVX1 U53 ( .A(a[8]), .Y(n27) );
  INVX1 U54 ( .A(n27), .Y(n28) );
  INVX1 U55 ( .A(n27), .Y(n29) );
  INVX1 U56 ( .A(a[9]), .Y(n30) );
  INVX1 U57 ( .A(n30), .Y(n31) );
  INVX1 U58 ( .A(n30), .Y(n32) );
  INVX1 U59 ( .A(a[10]), .Y(n33) );
  INVX1 U60 ( .A(n33), .Y(n34) );
  INVX1 U61 ( .A(n33), .Y(n35) );
  AND2X2 U62 ( .A(n34), .B(n14), .Y(n111) );
  INVX1 U63 ( .A(b[9]), .Y(n36) );
  INVX1 U64 ( .A(n36), .Y(n37) );
  INVX1 U65 ( .A(n36), .Y(n38) );
  INVX1 U66 ( .A(n321), .Y(n39) );
  NAND2BX1 U67 ( .AN(a[12]), .B(a[11]), .Y(n381) );
  BUFX3 U68 ( .A(n381), .Y(n92) );
  NAND2X1 U69 ( .A(b[0]), .B(n48), .Y(n47) );
  NAND2X1 U70 ( .A(b[0]), .B(n48), .Y(n63) );
  BUFX3 U71 ( .A(a[12]), .Y(n49) );
  NOR2BXL U72 ( .AN(a[12]), .B(n102), .Y(n108) );
  BUFX3 U73 ( .A(a[11]), .Y(n50) );
  INVX1 U74 ( .A(b[0]), .Y(n51) );
  NAND2X1 U75 ( .A(n34), .B(n102), .Y(n315) );
  XNOR3X2 U76 ( .A(n175), .B(n52), .C(n53), .Y(n265) );
  XNOR3X2 U77 ( .A(n163), .B(n229), .C(n82), .Y(n52) );
  XNOR3X2 U78 ( .A(n174), .B(n173), .C(n170), .Y(n53) );
  INVXL U79 ( .A(n376), .Y(n143) );
  NOR2XL U80 ( .A(n61), .B(n321), .Y(n323) );
  XOR2X1 U81 ( .A(n79), .B(n218), .Y(c[2]) );
  INVXL U82 ( .A(n102), .Y(n122) );
  OAI2BB1XL U83 ( .A0N(n50), .A1N(n122), .B0(n92), .Y(n128) );
  AOI22XL U84 ( .A0(n22), .A1(n199), .B0(n24), .B1(n200), .Y(n197) );
  AOI22XL U85 ( .A0(n29), .A1(n44), .B0(n32), .B1(n45), .Y(n42) );
  NAND2XL U86 ( .A(n100), .B(n107), .Y(n393) );
  AOI22XL U87 ( .A0(n35), .A1(n344), .B0(n32), .B1(n345), .Y(n342) );
  NAND2XL U88 ( .A(n97), .B(a[6]), .Y(n341) );
  NAND2XL U89 ( .A(b[8]), .B(n34), .Y(n236) );
  NAND2XL U90 ( .A(n38), .B(n35), .Y(n254) );
  NAND2XL U91 ( .A(n106), .B(n101), .Y(n229) );
  NAND2BXL U92 ( .AN(n95), .B(a[11]), .Y(n144) );
  NAND2XL U93 ( .A(n92), .B(n144), .Y(n147) );
  NAND2BXL U94 ( .AN(n99), .B(n49), .Y(n217) );
  NAND2XL U95 ( .A(n35), .B(n101), .Y(n54) );
  XNOR2X1 U96 ( .A(n297), .B(n296), .Y(n55) );
  NAND2XL U97 ( .A(n13), .B(n104), .Y(n152) );
  NAND2XL U98 ( .A(a[3]), .B(n102), .Y(n151) );
  NAND2XL U99 ( .A(n105), .B(n37), .Y(n391) );
  NAND2XL U100 ( .A(n106), .B(b[8]), .Y(n390) );
  NOR2X1 U101 ( .A(n234), .B(n233), .Y(n239) );
  AOI21XL U102 ( .A0(n92), .A1(n230), .B0(n389), .Y(n233) );
  NAND2XL U103 ( .A(a[7]), .B(n38), .Y(n208) );
  NAND2XL U104 ( .A(n49), .B(n14), .Y(n367) );
  NAND2XL U105 ( .A(n95), .B(n35), .Y(n287) );
  NAND2BXL U106 ( .AN(b[8]), .B(n50), .Y(n298) );
  NAND2XL U107 ( .A(n92), .B(n298), .Y(n301) );
  NAND2XL U108 ( .A(a[7]), .B(n19), .Y(n235) );
  NAND2XL U109 ( .A(n105), .B(n101), .Y(n256) );
  AOI22XL U110 ( .A0(n26), .A1(n75), .B0(n29), .B1(n76), .Y(n71) );
  NAND2XL U111 ( .A(n16), .B(n22), .Y(n81) );
  NAND2XL U112 ( .A(a[4]), .B(n10), .Y(n335) );
  NAND2XL U113 ( .A(n96), .B(n26), .Y(n340) );
  NAND2XL U114 ( .A(n107), .B(n39), .Y(n209) );
  NAND2XL U115 ( .A(a[3]), .B(n15), .Y(n89) );
  NAND2XL U116 ( .A(n99), .B(n35), .Y(n179) );
  NAND2XL U117 ( .A(b[8]), .B(n28), .Y(n180) );
  NAND2XL U118 ( .A(n100), .B(n31), .Y(n181) );
  NAND2XL U119 ( .A(n37), .B(n32), .Y(n237) );
  NAND2XL U120 ( .A(n38), .B(n319), .Y(n322) );
  NAND2XL U121 ( .A(n31), .B(n13), .Y(n316) );
  NAND2XL U122 ( .A(n15), .B(a[1]), .Y(n157) );
  INVXL U123 ( .A(n100), .Y(n389) );
  NAND2XL U124 ( .A(n106), .B(n14), .Y(n214) );
  NAND2XL U125 ( .A(n99), .B(n107), .Y(n294) );
  NAND2XL U126 ( .A(n106), .B(n37), .Y(n255) );
  NAND2XL U127 ( .A(a[7]), .B(n101), .Y(n171) );
  NAND2XL U128 ( .A(n104), .B(n97), .Y(n116) );
  NAND2XL U129 ( .A(n31), .B(n102), .Y(n296) );
  NAND2XL U130 ( .A(n29), .B(n19), .Y(n260) );
  NAND2XL U131 ( .A(n107), .B(n14), .Y(n225) );
  NAND2XL U132 ( .A(a[7]), .B(b[8]), .Y(n231) );
  NOR2BXL U133 ( .AN(n49), .B(n14), .Y(n126) );
  NAND2XL U134 ( .A(b[3]), .B(a[6]), .Y(n40) );
  NAND2XL U135 ( .A(n100), .B(n34), .Y(n215) );
  NAND2XL U136 ( .A(n29), .B(n101), .Y(n226) );
  NAND2XL U137 ( .A(n104), .B(b[3]), .Y(n156) );
  NAND2XL U138 ( .A(n107), .B(n102), .Y(n172) );
  NAND2XL U139 ( .A(n28), .B(n13), .Y(n297) );
  AND2X1 U140 ( .A(n96), .B(a[1]), .Y(n211) );
  INVXL U141 ( .A(n106), .Y(n387) );
  XNOR3X2 U142 ( .A(n57), .B(n58), .C(n221), .Y(n222) );
  NAND2XL U143 ( .A(n37), .B(n29), .Y(n57) );
  NAND2XL U144 ( .A(n18), .B(n32), .Y(n58) );
  NAND2XL U145 ( .A(n100), .B(a[7]), .Y(n257) );
  NAND2XL U146 ( .A(n99), .B(n26), .Y(n392) );
  NAND2BXL U147 ( .AN(n99), .B(n50), .Y(n230) );
  NAND2XL U148 ( .A(n100), .B(n24), .Y(n356) );
  NAND2XL U149 ( .A(n106), .B(n98), .Y(n355) );
  NAND2XL U150 ( .A(n96), .B(n32), .Y(n284) );
  NAND2XL U151 ( .A(n97), .B(n29), .Y(n285) );
  NAND2XL U152 ( .A(n98), .B(a[1]), .Y(n124) );
  NAND2XL U153 ( .A(n99), .B(n103), .Y(n125) );
  AOI22XL U154 ( .A0(n35), .A1(n312), .B0(n50), .B1(n313), .Y(n309) );
  NAND2XL U155 ( .A(b[3]), .B(n29), .Y(n307) );
  OAI2BB1XL U156 ( .A0N(n50), .A1N(n216), .B0(n92), .Y(n220) );
  XOR3X2 U157 ( .A(n59), .B(n303), .C(n361), .Y(n304) );
  NAND2XL U158 ( .A(n16), .B(n21), .Y(n59) );
  NAND2XL U159 ( .A(a[0]), .B(n14), .Y(n279) );
  AOI22XL U160 ( .A0(a[6]), .A1(n93), .B0(n26), .B1(n94), .Y(n90) );
  NAND2XL U161 ( .A(n105), .B(b[3]), .Y(n88) );
  INVXL U162 ( .A(n96), .Y(n394) );
  XOR3X2 U163 ( .A(n60), .B(n354), .C(n353), .Y(n358) );
  NAND2XL U164 ( .A(n29), .B(n95), .Y(n60) );
  NAND2XL U165 ( .A(n14), .B(a[1]), .Y(n136) );
  NAND2XL U166 ( .A(n102), .B(n104), .Y(n137) );
  NAND2XL U167 ( .A(n101), .B(a[3]), .Y(n138) );
  NOR2BXL U168 ( .AN(n50), .B(n97), .Y(n189) );
  NAND2XL U169 ( .A(n99), .B(n28), .Y(n85) );
  NAND2XL U170 ( .A(n31), .B(n98), .Y(n86) );
  NAND2XL U171 ( .A(n28), .B(n98), .Y(n83) );
  NAND2XL U172 ( .A(n32), .B(n97), .Y(n84) );
  NAND2XL U173 ( .A(n18), .B(n21), .Y(n347) );
  NAND2XL U174 ( .A(a[3]), .B(n96), .Y(n115) );
  NAND2XL U175 ( .A(n98), .B(n26), .Y(n293) );
  XOR2X1 U176 ( .A(n263), .B(n262), .Y(n291) );
  NAND2XL U177 ( .A(n26), .B(n14), .Y(n261) );
  AOI22XL U178 ( .A0(n24), .A1(n185), .B0(n105), .B1(n186), .Y(n183) );
  NAND2XL U179 ( .A(a[5]), .B(b[3]), .Y(n69) );
  NAND2XL U180 ( .A(n105), .B(n14), .Y(n207) );
  NAND2XL U181 ( .A(n106), .B(n102), .Y(n206) );
  NAND2XL U182 ( .A(n103), .B(n19), .Y(n368) );
  INVXL U183 ( .A(n98), .Y(n216) );
  AND2X1 U184 ( .A(n105), .B(n102), .Y(n82) );
  AND2X1 U185 ( .A(n35), .B(n97), .Y(n150) );
  AND2X1 U186 ( .A(n35), .B(n96), .Y(n135) );
  AND2X1 U187 ( .A(n32), .B(n101), .Y(n259) );
  AND2X1 U188 ( .A(n103), .B(n97), .Y(n212) );
  AND2X1 U189 ( .A(n103), .B(n18), .Y(n329) );
  AND2X1 U190 ( .A(n26), .B(n95), .Y(n43) );
  INVXL U191 ( .A(n50), .Y(n378) );
  AND2X1 U192 ( .A(n92), .B(n318), .Y(n61) );
  NAND2XL U193 ( .A(n11), .B(n104), .Y(n339) );
  NAND2XL U194 ( .A(n105), .B(n15), .Y(n70) );
  INVXL U195 ( .A(n107), .Y(n74) );
  NAND2XL U196 ( .A(n16), .B(n24), .Y(n338) );
  NAND2XL U197 ( .A(a[6]), .B(n10), .Y(n364) );
  NAND2XL U198 ( .A(a[5]), .B(n16), .Y(n365) );
  NAND2XL U199 ( .A(a[4]), .B(n11), .Y(n366) );
  NAND2XL U200 ( .A(n15), .B(n26), .Y(n308) );
  NAND2XL U201 ( .A(n103), .B(n38), .Y(n343) );
  NAND2XL U202 ( .A(n24), .B(n18), .Y(n328) );
  NAND2XL U203 ( .A(n15), .B(a[5]), .Y(n41) );
  NAND2XL U204 ( .A(a[4]), .B(n16), .Y(n351) );
  NAND2XL U205 ( .A(n103), .B(n11), .Y(n289) );
  NAND2XL U206 ( .A(n24), .B(n95), .Y(n158) );
  NAND2XL U207 ( .A(n18), .B(n104), .Y(n352) );
  NAND2XL U208 ( .A(n103), .B(n10), .Y(n246) );
  NAND2XL U209 ( .A(n10), .B(n24), .Y(n311) );
  NAND2XL U210 ( .A(n11), .B(n21), .Y(n306) );
  NAND2XL U211 ( .A(n22), .B(n39), .Y(n273) );
  NAND2XL U212 ( .A(n21), .B(n19), .Y(n274) );
  NAND2XL U213 ( .A(a[4]), .B(n18), .Y(n275) );
  NAND2XL U214 ( .A(n24), .B(n38), .Y(n276) );
  AND2X1 U215 ( .A(n21), .B(n39), .Y(n87) );
  NAND2BXL U216 ( .AN(b[1]), .B(n50), .Y(n129) );
  NAND2XL U217 ( .A(n92), .B(n129), .Y(n132) );
  INVXL U218 ( .A(b[1]), .Y(n380) );
  NAND2X1 U219 ( .A(b[1]), .B(n46), .Y(n62) );
  XNOR2X1 U220 ( .A(n143), .B(n176), .Y(n360) );
  XNOR2X1 U221 ( .A(n68), .B(n8), .Y(n314) );
  XOR2X1 U222 ( .A(n143), .B(n377), .Y(n64) );
  XOR3X2 U223 ( .A(n361), .B(n360), .C(n359), .Y(c[10]) );
  NAND3X1 U224 ( .A(n61), .B(n320), .C(n322), .Y(n326) );
  XOR2X1 U225 ( .A(n232), .B(n231), .Y(n175) );
  XNOR3X2 U226 ( .A(n64), .B(n177), .C(n203), .Y(n223) );
  XNOR3X2 U227 ( .A(n334), .B(n333), .C(n332), .Y(c[8]) );
  XOR3X2 U228 ( .A(n204), .B(n264), .C(n203), .Y(n205) );
  XNOR3X2 U229 ( .A(n314), .B(n79), .C(n249), .Y(c[5]) );
  XNOR3X2 U230 ( .A(n159), .B(n248), .C(n247), .Y(n249) );
  XOR2X1 U231 ( .A(n246), .B(n158), .Y(n247) );
  XNOR2X1 U232 ( .A(n156), .B(n157), .Y(n248) );
  INVX1 U233 ( .A(n367), .Y(n377) );
  NOR2X1 U234 ( .A(n387), .B(n389), .Y(n295) );
  XOR3X2 U235 ( .A(n65), .B(n66), .C(n67), .Y(n359) );
  XNOR3X2 U236 ( .A(n340), .B(n341), .C(n342), .Y(n65) );
  XOR2X1 U237 ( .A(n352), .B(n351), .Y(n66) );
  XNOR2X1 U238 ( .A(n358), .B(n357), .Y(n67) );
  INVX1 U239 ( .A(n370), .Y(n176) );
  XOR2X1 U240 ( .A(n226), .B(n225), .Y(n240) );
  XOR3X2 U241 ( .A(n237), .B(n236), .C(n235), .Y(n238) );
  XNOR3X2 U242 ( .A(n377), .B(n265), .C(n264), .Y(n266) );
  XOR3X2 U243 ( .A(n77), .B(n78), .C(n222), .Y(n68) );
  XNOR2X1 U244 ( .A(n215), .B(n214), .Y(n77) );
  XOR2X1 U245 ( .A(n172), .B(n171), .Y(n78) );
  XNOR3X2 U246 ( .A(n80), .B(n278), .C(n266), .Y(c[6]) );
  XOR2X1 U247 ( .A(n112), .B(n123), .Y(n278) );
  XOR2X1 U248 ( .A(n269), .B(n270), .Y(c[12]) );
  XOR2X1 U249 ( .A(n271), .B(n272), .Y(n270) );
  XOR2X1 U250 ( .A(n372), .B(n371), .Y(n373) );
  XNOR3X2 U251 ( .A(n328), .B(n7), .C(n369), .Y(n372) );
  XOR3X2 U252 ( .A(n308), .B(n370), .C(n87), .Y(n371) );
  INVX1 U253 ( .A(n381), .Y(n188) );
  XNOR2X1 U254 ( .A(n291), .B(n8), .Y(n80) );
  XOR2XL U255 ( .A(n291), .B(n6), .Y(n361) );
  XOR2X1 U256 ( .A(n305), .B(n304), .Y(c[7]) );
  XOR2X1 U257 ( .A(n210), .B(n205), .Y(c[3]) );
  XNOR3X2 U258 ( .A(n80), .B(n350), .C(n349), .Y(c[9]) );
  XOR3X2 U259 ( .A(n375), .B(n374), .C(n373), .Y(c[11]) );
  NOR2XL U260 ( .A(n73), .B(n387), .Y(n91) );
  OAI21XL U261 ( .A0(n32), .A1(n380), .B0(n9), .Y(n44) );
  OAI21XL U262 ( .A0(n29), .A1(n46), .B0(n47), .Y(n45) );
  OAI21XL U263 ( .A0(n24), .A1(n48), .B0(n9), .Y(n199) );
  OAI21XL U264 ( .A0(n104), .A1(n51), .B0(n47), .Y(n200) );
  AOI22X1 U265 ( .A0(n106), .A1(n120), .B0(n107), .B1(n121), .Y(n117) );
  OAI21XL U266 ( .A0(n107), .A1(n380), .B0(n9), .Y(n120) );
  OAI21XL U267 ( .A0(n106), .A1(n46), .B0(n63), .Y(n121) );
  OAI21XL U268 ( .A0(n35), .A1(n380), .B0(n62), .Y(n345) );
  OAI21XL U269 ( .A0(n32), .A1(n51), .B0(n47), .Y(n344) );
  OAI2BB1X1 U270 ( .A0N(n14), .A1N(n128), .B0(n127), .Y(n370) );
  INVXL U271 ( .A(n99), .Y(n227) );
  XOR2X2 U272 ( .A(n202), .B(n196), .Y(n264) );
  XNOR3X2 U273 ( .A(n209), .B(n208), .C(n195), .Y(n196) );
  NAND3X1 U274 ( .A(n194), .B(n193), .C(n192), .Y(n202) );
  OAI21XL U275 ( .A0(n21), .A1(n51), .B0(n47), .Y(n244) );
  OAI21XL U276 ( .A0(n24), .A1(n51), .B0(n47), .Y(n186) );
  OAI21XL U277 ( .A0(n26), .A1(n51), .B0(n47), .Y(n76) );
  OAI21XL U278 ( .A0(n106), .A1(n48), .B0(n9), .Y(n160) );
  OAI21XL U279 ( .A0(n105), .A1(n51), .B0(n47), .Y(n161) );
  OAI21XL U280 ( .A0(a[6]), .A1(n51), .B0(n47), .Y(n94) );
  OAI21XL U281 ( .A0(n35), .A1(n51), .B0(n47), .Y(n313) );
  OAI2BB1X2 U282 ( .A0N(n102), .A1N(n110), .B0(n109), .Y(n119) );
  OAI21XL U283 ( .A0(n105), .A1(n48), .B0(n62), .Y(n185) );
  OAI21XL U284 ( .A0(n29), .A1(n380), .B0(n9), .Y(n75) );
  OAI21XL U285 ( .A0(n50), .A1(n48), .B0(n62), .Y(n312) );
  XNOR3X2 U286 ( .A(n256), .B(n154), .C(n153), .Y(n155) );
  XNOR3X2 U287 ( .A(n150), .B(n149), .C(n148), .Y(n162) );
  INVX1 U288 ( .A(n95), .Y(n73) );
  OAI2BB1X1 U289 ( .A0N(n96), .A1N(n147), .B0(n146), .Y(n149) );
  XOR2X1 U290 ( .A(n261), .B(n260), .Y(n262) );
  XNOR3X2 U291 ( .A(n259), .B(n254), .C(n253), .Y(n263) );
  NOR2BX1 U292 ( .AN(a[11]), .B(n96), .Y(n167) );
  XNOR2X1 U293 ( .A(n316), .B(n315), .Y(n324) );
  XOR2X1 U294 ( .A(n142), .B(n141), .Y(n203) );
  XNOR3X2 U295 ( .A(n393), .B(n140), .C(n139), .Y(n141) );
  XNOR3X2 U296 ( .A(n135), .B(n134), .C(n133), .Y(n142) );
  XNOR3X2 U297 ( .A(n376), .B(n337), .C(n336), .Y(n350) );
  XOR2X1 U298 ( .A(n335), .B(n41), .Y(n336) );
  XNOR2X1 U299 ( .A(n40), .B(n43), .Y(n337) );
  NOR2BX1 U300 ( .AN(n49), .B(n98), .Y(n182) );
  XNOR3X2 U301 ( .A(n81), .B(n71), .C(n314), .Y(n333) );
  XOR2X1 U302 ( .A(n290), .B(n289), .Y(n303) );
  NAND2X1 U303 ( .A(n98), .B(n104), .Y(n290) );
  XNOR3X2 U304 ( .A(n224), .B(n286), .C(n223), .Y(c[4]) );
  XOR2X1 U305 ( .A(n183), .B(n213), .Y(n224) );
  XOR3X2 U306 ( .A(n212), .B(n211), .C(n184), .Y(n213) );
  OAI2BB1X1 U307 ( .A0N(n38), .A1N(n301), .B0(n300), .Y(n302) );
  XOR2X1 U308 ( .A(n165), .B(n164), .Y(n173) );
  NAND2X1 U309 ( .A(n100), .B(n28), .Y(n165) );
  NAND2X1 U310 ( .A(n99), .B(n31), .Y(n164) );
  XOR2X1 U311 ( .A(n152), .B(n151), .Y(n154) );
  XOR2X1 U312 ( .A(n391), .B(n390), .Y(n140) );
  XOR3X2 U313 ( .A(n279), .B(n277), .C(n386), .Y(n269) );
  XOR2X1 U314 ( .A(n280), .B(n281), .Y(n277) );
  XOR2X1 U315 ( .A(n282), .B(n283), .Y(n281) );
  XNOR3X2 U316 ( .A(n90), .B(n288), .C(n286), .Y(n305) );
  XOR3X2 U317 ( .A(n89), .B(n88), .C(n91), .Y(n288) );
  XNOR3X2 U318 ( .A(n64), .B(n201), .C(n178), .Y(n210) );
  NOR2X1 U319 ( .A(n388), .B(n394), .Y(n201) );
  XNOR2X1 U320 ( .A(n198), .B(n197), .Y(n178) );
  XOR2X1 U321 ( .A(n284), .B(n285), .Y(n283) );
  NAND2X1 U322 ( .A(n107), .B(n37), .Y(n232) );
  XNOR3X2 U323 ( .A(n309), .B(n363), .C(n362), .Y(n375) );
  XNOR2X1 U324 ( .A(n310), .B(n307), .Y(n362) );
  OAI2BB1X1 U325 ( .A0N(n96), .A1N(n169), .B0(n168), .Y(n170) );
  OAI21XL U326 ( .A0(n167), .A1(n188), .B0(n97), .Y(n168) );
  INVX1 U327 ( .A(n97), .Y(n166) );
  NAND2BX1 U328 ( .AN(n63), .B(n49), .Y(n384) );
  XNOR3X2 U329 ( .A(n83), .B(n84), .C(n392), .Y(n133) );
  XOR3X2 U330 ( .A(n138), .B(n137), .C(n136), .Y(n139) );
  XOR2X1 U331 ( .A(n241), .B(n242), .Y(n218) );
  NOR2X1 U332 ( .A(n388), .B(n73), .Y(n242) );
  AOI22X1 U333 ( .A0(n21), .A1(n243), .B0(n22), .B1(n244), .Y(n241) );
  OAI21XL U334 ( .A0(n22), .A1(n380), .B0(n62), .Y(n243) );
  OAI2BB1X1 U335 ( .A0N(n18), .A1N(n252), .B0(n251), .Y(n253) );
  AOI21X1 U336 ( .A0(n99), .A1(n220), .B0(n219), .Y(n221) );
  XOR3X2 U337 ( .A(n181), .B(n180), .C(n179), .Y(n191) );
  XNOR3X2 U338 ( .A(n379), .B(n360), .C(n203), .Y(c[0]) );
  NOR2X1 U339 ( .A(n388), .B(n51), .Y(n379) );
  XOR2X1 U340 ( .A(n385), .B(n287), .Y(n282) );
  XOR2X1 U341 ( .A(n395), .B(n292), .Y(n280) );
  XOR2X1 U342 ( .A(n293), .B(n294), .Y(n292) );
  XOR3X2 U343 ( .A(n295), .B(n377), .C(n376), .Y(n395) );
  XOR2X1 U344 ( .A(n113), .B(n114), .Y(n112) );
  XOR2X1 U345 ( .A(n115), .B(n116), .Y(n114) );
  XOR2X1 U346 ( .A(n117), .B(n118), .Y(n113) );
  NOR2BX1 U347 ( .AN(n49), .B(n38), .Y(n299) );
  NOR2BX1 U348 ( .AN(a[12]), .B(n96), .Y(n145) );
  OAI21XL U349 ( .A0(n189), .A1(n188), .B0(n98), .Y(n190) );
  NOR2BX1 U350 ( .AN(n49), .B(n18), .Y(n250) );
  NOR2BX1 U351 ( .AN(n49), .B(n95), .Y(n130) );
  XNOR3X2 U352 ( .A(n348), .B(n347), .C(n346), .Y(n349) );
  XOR3X2 U353 ( .A(n343), .B(n339), .C(n338), .Y(n346) );
  XOR2X1 U354 ( .A(n386), .B(n42), .Y(n348) );
  NAND2BXL U355 ( .AN(n100), .B(n49), .Y(n228) );
  AND2X2 U356 ( .A(n13), .B(a[3]), .Y(n163) );
  XNOR3X2 U357 ( .A(n85), .B(n86), .C(n257), .Y(n148) );
  AND2X2 U358 ( .A(n34), .B(n98), .Y(n174) );
  NAND2BXL U359 ( .AN(n37), .B(a[11]), .Y(n318) );
  XNOR2X1 U360 ( .A(n255), .B(n258), .Y(n153) );
  XNOR2X1 U361 ( .A(n207), .B(n206), .Y(n195) );
  XNOR2X1 U362 ( .A(n331), .B(n330), .Y(n332) );
  XOR2X1 U363 ( .A(n69), .B(n72), .Y(n330) );
  XNOR3X2 U364 ( .A(n329), .B(n70), .C(n363), .Y(n331) );
  INVX1 U365 ( .A(n101), .Y(n321) );
  OAI21XL U366 ( .A0(n26), .A1(n380), .B0(n62), .Y(n93) );
  NOR2X1 U367 ( .A(n73), .B(n74), .Y(n72) );
  NOR2X1 U368 ( .A(n73), .B(n56), .Y(n184) );
  INVX1 U369 ( .A(n104), .Y(n56) );
  XOR2X1 U370 ( .A(n311), .B(n306), .Y(n334) );
  NOR2BX1 U371 ( .AN(n32), .B(n73), .Y(n310) );
  XNOR3X2 U372 ( .A(n366), .B(n365), .C(n364), .Y(n374) );
  NAND2X1 U373 ( .A(n38), .B(a[1]), .Y(n353) );
  NAND2X1 U374 ( .A(n103), .B(n39), .Y(n354) );
  XOR2X1 U375 ( .A(n356), .B(n355), .Y(n357) );
  XOR2X1 U376 ( .A(n273), .B(n274), .Y(n272) );
  XOR2X1 U377 ( .A(n124), .B(n125), .Y(n123) );
  INVX1 U378 ( .A(n103), .Y(n388) );
  XOR2X1 U379 ( .A(n275), .B(n276), .Y(n271) );
  AOI22X1 U380 ( .A0(a[0]), .A1(n267), .B0(n21), .B1(n268), .Y(n245) );
  OAI21XL U381 ( .A0(n21), .A1(n48), .B0(n9), .Y(n267) );
  OAI21XL U382 ( .A0(n103), .A1(n51), .B0(n47), .Y(n268) );
  XOR2X1 U383 ( .A(n368), .B(n367), .Y(n369) );
  INVX1 U384 ( .A(b[0]), .Y(n46) );
  OAI2BB1X1 U385 ( .A0N(n95), .A1N(n132), .B0(n131), .Y(n134) );
  BUFX3 U386 ( .A(a[4]), .Y(n105) );
  BUFX3 U387 ( .A(a[6]), .Y(n107) );
  BUFX3 U388 ( .A(a[2]), .Y(n104) );
  BUFX3 U389 ( .A(a[5]), .Y(n106) );
  BUFX3 U390 ( .A(b[10]), .Y(n101) );
  BUFX3 U391 ( .A(b[11]), .Y(n102) );
  BUFX3 U392 ( .A(b[3]), .Y(n96) );
  BUFX3 U393 ( .A(b[4]), .Y(n97) );
  BUFX3 U394 ( .A(b[5]), .Y(n98) );
  BUFX3 U395 ( .A(b[6]), .Y(n99) );
  BUFX3 U396 ( .A(b[7]), .Y(n100) );
  INVX1 U397 ( .A(b[1]), .Y(n48) );
  BUFX3 U398 ( .A(a[0]), .Y(n103) );
  BUFX3 U399 ( .A(b[2]), .Y(n95) );
  OAI21XL U400 ( .A0(n126), .A1(n382), .B0(n19), .Y(n127) );
  OAI21XL U401 ( .A0(n182), .A1(n382), .B0(n97), .Y(n187) );
  OAI21XL U402 ( .A0(n299), .A1(n382), .B0(n18), .Y(n300) );
  AOI21XL U403 ( .A0(n317), .A1(n217), .B0(n216), .Y(n219) );
  OAI21XL U404 ( .A0(n130), .A1(n382), .B0(b[1]), .Y(n131) );
  AOI21XL U405 ( .A0(n317), .A1(n228), .B0(n227), .Y(n234) );
  OAI21XL U406 ( .A0(n250), .A1(n382), .B0(n100), .Y(n251) );
  AOI2BB2X1 U407 ( .B0(b[0]), .B1(n382), .A0N(n92), .A1N(n380), .Y(n383) );
  OAI2BB1XL U408 ( .A0N(a[12]), .A1N(n166), .B0(n317), .Y(n169) );
endmodule


module degree_computation_3 ( deg_Ri, deg_Qi, stop_i, d1out, start, deg_Ro, 
        deg_Qo, stop_o, sw, clk, reset );
  input [4:0] deg_Ri;
  input [4:0] deg_Qi;
  input [12:0] d1out;
  output [4:0] deg_Ro;
  output [4:0] deg_Qo;
  input stop_i, start, clk, reset;
  output stop_o, sw;
  wire   out, sw_reg, stop2_signal, n2, n3, n4, n5, n6, n1, n7, n8, n9, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22;
  wire   [4:0] DQ1;
  wire   [4:0] DR1;
  wire   [4:0] rmux_signal;
  wire   [4:0] qmux_signal;
  wire   [4:0] DR2;
  wire   [4:0] addr_signal;
  wire   [4:0] DQ2;
  wire   [4:0] addq_signal;
  wire   [4:0] mr_signal;
  wire   [4:0] mq_signal;
  wire   [4:0] r2mux_signal;
  wire   [4:0] q2mux_signal;
  wire   [12:0] dmux_signal;

  mux_5_23 mdeg1 ( .a(DQ1), .b(DR1), .sel(sw_reg), .out(rmux_signal) );
  mux_5_22 mdeg2 ( .a(DR1), .b(DQ1), .sel(n9), .out(qmux_signal) );
  mux_5_21 mdeg3 ( .a(DR2), .b(addr_signal), .sel(n8), .out(mr_signal) );
  mux_5_20 mdeg4 ( .a(addq_signal), .b(DQ2), .sel(n7), .out(mq_signal) );
  mux_5_19 mdeg5 ( .a(DR2), .b(mr_signal), .sel(n11), .out(r2mux_signal) );
  mux_5_18 mdeg6 ( .a(DQ2), .b(mq_signal), .sel(n11), .out(q2mux_signal) );
  mux_13_19 mdeg7 ( .a(d1out), .b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .sel(stop2_signal), .out(
        dmux_signal) );
  degree_computation_3_DW01_dec_0 sub_41 ( .A(DQ2), .SUM(addq_signal) );
  degree_computation_3_DW01_dec_1 sub_40 ( .A(DR2), .SUM(addr_signal) );
  DFFRHQX1 \DQ3_reg[2]  ( .D(q2mux_signal[2]), .CK(clk), .RN(reset), .Q(
        deg_Qo[2]) );
  DFFRHQX1 \DQ3_reg[3]  ( .D(q2mux_signal[3]), .CK(clk), .RN(reset), .Q(
        deg_Qo[3]) );
  DFFRHQX1 \DQ3_reg[4]  ( .D(q2mux_signal[4]), .CK(clk), .RN(reset), .Q(
        deg_Qo[4]) );
  DFFRHQX1 \DR3_reg[1]  ( .D(r2mux_signal[1]), .CK(clk), .RN(reset), .Q(
        deg_Ro[1]) );
  DFFRHQX1 \DR3_reg[0]  ( .D(r2mux_signal[0]), .CK(clk), .RN(reset), .Q(
        deg_Ro[0]) );
  DFFRHQX1 \DQ3_reg[0]  ( .D(q2mux_signal[0]), .CK(clk), .RN(reset), .Q(
        deg_Qo[0]) );
  DFFRHQX1 \DR3_reg[3]  ( .D(r2mux_signal[3]), .CK(clk), .RN(reset), .Q(
        deg_Ro[3]) );
  DFFRHQX1 \DR3_reg[4]  ( .D(r2mux_signal[4]), .CK(clk), .RN(reset), .Q(
        deg_Ro[4]) );
  DFFRHQX1 \DQ3_reg[1]  ( .D(q2mux_signal[1]), .CK(clk), .RN(reset), .Q(
        deg_Qo[1]) );
  DFFRHQX1 \DR3_reg[2]  ( .D(r2mux_signal[2]), .CK(clk), .RN(reset), .Q(
        deg_Ro[2]) );
  DFFRHQX1 \DQ1_reg[3]  ( .D(deg_Qi[3]), .CK(clk), .RN(reset), .Q(DQ1[3]) );
  DFFRHQX1 \DQ1_reg[2]  ( .D(deg_Qi[2]), .CK(clk), .RN(reset), .Q(DQ1[2]) );
  DFFRHQX1 \DQ1_reg[1]  ( .D(deg_Qi[1]), .CK(clk), .RN(reset), .Q(DQ1[1]) );
  DFFRHQX1 \DQ1_reg[0]  ( .D(deg_Qi[0]), .CK(clk), .RN(reset), .Q(DQ1[0]) );
  DFFRHQX1 \DR1_reg[3]  ( .D(deg_Ri[3]), .CK(clk), .RN(reset), .Q(DR1[3]) );
  DFFRHQX1 \DR1_reg[2]  ( .D(deg_Ri[2]), .CK(clk), .RN(reset), .Q(DR1[2]) );
  DFFRHQX1 \DR1_reg[1]  ( .D(deg_Ri[1]), .CK(clk), .RN(reset), .Q(DR1[1]) );
  DFFRHQX1 \DR1_reg[0]  ( .D(deg_Ri[0]), .CK(clk), .RN(reset), .Q(DR1[0]) );
  DFFRHQX1 \DQ1_reg[4]  ( .D(deg_Qi[4]), .CK(clk), .RN(reset), .Q(DQ1[4]) );
  DFFRHQX1 \DR1_reg[4]  ( .D(deg_Ri[4]), .CK(clk), .RN(reset), .Q(DR1[4]) );
  DFFRHQX1 \DQ2_reg[4]  ( .D(qmux_signal[4]), .CK(clk), .RN(reset), .Q(DQ2[4])
         );
  DFFRHQX1 \DR2_reg[4]  ( .D(rmux_signal[4]), .CK(clk), .RN(reset), .Q(DR2[4])
         );
  DFFRHQX1 sw_reg_reg ( .D(out), .CK(clk), .RN(reset), .Q(sw_reg) );
  DFFRHQX1 shift_reg_reg ( .D(out), .CK(clk), .RN(reset), .Q(sw) );
  DFFRHQX1 \DQ2_reg[2]  ( .D(qmux_signal[2]), .CK(clk), .RN(reset), .Q(DQ2[2])
         );
  DFFRHQX1 \DR2_reg[2]  ( .D(rmux_signal[2]), .CK(clk), .RN(reset), .Q(DR2[2])
         );
  DFFRHQX1 \DQ2_reg[1]  ( .D(qmux_signal[1]), .CK(clk), .RN(reset), .Q(DQ2[1])
         );
  DFFRHQX1 \DR2_reg[1]  ( .D(rmux_signal[1]), .CK(clk), .RN(reset), .Q(DR2[1])
         );
  DFFRHQX1 \DQ2_reg[3]  ( .D(qmux_signal[3]), .CK(clk), .RN(reset), .Q(DQ2[3])
         );
  DFFRHQX1 \DR2_reg[3]  ( .D(rmux_signal[3]), .CK(clk), .RN(reset), .Q(DR2[3])
         );
  DFFRHQX1 \DQ2_reg[0]  ( .D(qmux_signal[0]), .CK(clk), .RN(reset), .Q(DQ2[0])
         );
  DFFRHQX1 \DR2_reg[0]  ( .D(rmux_signal[0]), .CK(clk), .RN(reset), .Q(DR2[0])
         );
  DFFSX1 start_reg_reg ( .D(start), .CK(clk), .SN(reset), .Q(stop2_signal) );
  NAND4X1 U3 ( .A(n3), .B(n4), .C(n5), .D(n6), .Y(n1) );
  INVX1 U4 ( .A(n1), .Y(n7) );
  INVX1 U5 ( .A(n1), .Y(n8) );
  BUFX3 U6 ( .A(sw_reg), .Y(n9) );
  INVX1 U7 ( .A(n12), .Y(n11) );
  INVX1 U8 ( .A(stop_i), .Y(n12) );
  NOR3X1 U9 ( .A(dmux_signal[0]), .B(dmux_signal[11]), .C(dmux_signal[10]), 
        .Y(n3) );
  NOR3X1 U10 ( .A(dmux_signal[12]), .B(dmux_signal[2]), .C(dmux_signal[1]), 
        .Y(n4) );
  NOR3X1 U11 ( .A(dmux_signal[3]), .B(dmux_signal[5]), .C(dmux_signal[4]), .Y(
        n5) );
  NOR4X1 U12 ( .A(dmux_signal[9]), .B(dmux_signal[8]), .C(dmux_signal[7]), .D(
        dmux_signal[6]), .Y(n6) );
  AND2X2 U13 ( .A(stop2_signal), .B(n2), .Y(stop_o) );
  OAI22X1 U14 ( .A0(mr_signal[4]), .A1(mr_signal[3]), .B0(mq_signal[4]), .B1(
        mq_signal[3]), .Y(n2) );
  INVX1 U15 ( .A(deg_Qi[4]), .Y(n22) );
  INVX1 U16 ( .A(deg_Ri[1]), .Y(n15) );
  AOI2BB1X1 U17 ( .A0N(n15), .A1N(deg_Qi[1]), .B0(deg_Ri[0]), .Y(n14) );
  INVX1 U18 ( .A(deg_Qi[2]), .Y(n17) );
  INVX1 U19 ( .A(deg_Qi[3]), .Y(n13) );
  AND2X1 U20 ( .A(deg_Ri[3]), .B(n13), .Y(n16) );
  OAI32X1 U21 ( .A0(n17), .A1(deg_Ri[2]), .A2(n16), .B0(deg_Ri[3]), .B1(n13), 
        .Y(n18) );
  AOI221X1 U22 ( .A0(deg_Qi[1]), .A1(n15), .B0(n14), .B1(deg_Qi[0]), .C0(n18), 
        .Y(n21) );
  AOI21X1 U23 ( .A0(deg_Ri[2]), .A1(n17), .B0(n16), .Y(n19) );
  OAI2BB2X1 U24 ( .B0(n19), .B1(n18), .A0N(n22), .A1N(deg_Ri[4]), .Y(n20) );
  OAI22X1 U25 ( .A0(deg_Ri[4]), .A1(n22), .B0(n21), .B1(n20), .Y(out) );
endmodule


module multiplier_column8_p16 ( b, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, 
        P11, P12, P13, P14, P15, P16 );
  input [12:0] b;
  output [12:0] P1;
  output [12:0] P2;
  output [12:0] P3;
  output [12:0] P4;
  output [12:0] P5;
  output [12:0] P6;
  output [12:0] P7;
  output [12:0] P8;
  output [12:0] P9;
  output [12:0] P10;
  output [12:0] P11;
  output [12:0] P12;
  output [12:0] P13;
  output [12:0] P14;
  output [12:0] P15;
  output [12:0] P16;
  wire   b_3, b_2, b_1, b_0, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n37, n38, n39, n40,
         n41, n42, n43, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n157, n160, n1,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n35, n36, n44, n58,
         n110, n132, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199;
  assign b_3 = b[3];
  assign b_2 = b[2];
  assign b_1 = b[1];
  assign b_0 = b[0];

  XNOR2X4 U257 ( .A(n17), .B(b[9]), .Y(n51) );
  INVX2 U1 ( .A(n192), .Y(n94) );
  XNOR2X1 U2 ( .A(n94), .B(n189), .Y(n30) );
  XOR2X1 U3 ( .A(n190), .B(P12[11]), .Y(n109) );
  XOR2X1 U4 ( .A(n198), .B(n22), .Y(P9[11]) );
  XOR2XL U5 ( .A(n45), .B(P5[1]), .Y(P7[6]) );
  XNOR2X2 U6 ( .A(n20), .B(P10[3]), .Y(P14[9]) );
  XNOR2X2 U7 ( .A(P4[1]), .B(n13), .Y(P10[3]) );
  XNOR2X1 U8 ( .A(n126), .B(n94), .Y(n131) );
  INVX2 U9 ( .A(b[11]), .Y(n132) );
  BUFX3 U10 ( .A(b[11]), .Y(n197) );
  XNOR2X1 U11 ( .A(n94), .B(n191), .Y(n160) );
  XNOR2X4 U12 ( .A(n132), .B(b_1), .Y(n15) );
  XNOR2X1 U13 ( .A(n24), .B(n27), .Y(n118) );
  XNOR2X1 U14 ( .A(n6), .B(n15), .Y(n155) );
  XNOR2X1 U15 ( .A(P11[9]), .B(n193), .Y(n126) );
  XOR2X1 U16 ( .A(n4), .B(n155), .Y(P11[9]) );
  XOR2X1 U17 ( .A(n193), .B(n149), .Y(n34) );
  XOR2X1 U18 ( .A(n4), .B(n98), .Y(P12[5]) );
  XOR2X1 U19 ( .A(n188), .B(n150), .Y(P9[0]) );
  INVX1 U20 ( .A(b_0), .Y(n6) );
  INVX1 U21 ( .A(n187), .Y(n5) );
  BUFX3 U22 ( .A(b_0), .Y(n187) );
  CLKBUFX1 U23 ( .A(P16[0]), .Y(P15[5]) );
  INVX1 U24 ( .A(b[8]), .Y(n1) );
  BUFX4 U25 ( .A(b[8]), .Y(n195) );
  INVX1 U26 ( .A(n195), .Y(n42) );
  XNOR2XL U27 ( .A(n28), .B(n45), .Y(P11[8]) );
  BUFX3 U28 ( .A(b_1), .Y(n188) );
  INVX1 U29 ( .A(n94), .Y(P1[0]) );
  XOR2X1 U30 ( .A(n192), .B(n197), .Y(n116) );
  BUFX3 U31 ( .A(b[5]), .Y(n192) );
  XNOR2XL U32 ( .A(n193), .B(n78), .Y(P16[11]) );
  INVX1 U33 ( .A(n32), .Y(P1[12]) );
  BUFX3 U34 ( .A(b[12]), .Y(n4) );
  INVX4 U35 ( .A(n198), .Y(n17) );
  INVX1 U36 ( .A(n194), .Y(n7) );
  XNOR2XL U37 ( .A(n53), .B(n193), .Y(P1[2]) );
  INVX1 U38 ( .A(n194), .Y(n53) );
  INVX1 U39 ( .A(n189), .Y(n8) );
  INVX1 U40 ( .A(b[6]), .Y(n9) );
  INVXL U41 ( .A(n193), .Y(n10) );
  XNOR2X1 U42 ( .A(n187), .B(n10), .Y(n123) );
  XNOR2X1 U43 ( .A(n50), .B(n10), .Y(n70) );
  INVX1 U44 ( .A(b[9]), .Y(n11) );
  INVX1 U45 ( .A(b_3), .Y(n13) );
  INVX1 U46 ( .A(b_3), .Y(n12) );
  XNOR2XL U47 ( .A(n13), .B(n34), .Y(P2[9]) );
  XNOR2XL U48 ( .A(n12), .B(n41), .Y(P8[10]) );
  XNOR2X2 U49 ( .A(n65), .B(n12), .Y(n64) );
  XNOR2XL U50 ( .A(n12), .B(n192), .Y(n77) );
  XNOR2XL U51 ( .A(n13), .B(n155), .Y(n97) );
  XOR2XL U52 ( .A(n80), .B(n76), .Y(n100) );
  XNOR2X1 U53 ( .A(n112), .B(n189), .Y(n72) );
  XNOR2XL U54 ( .A(n189), .B(n9), .Y(n47) );
  XNOR2XL U55 ( .A(n4), .B(n193), .Y(n119) );
  BUFX3 U56 ( .A(b[12]), .Y(n198) );
  XNOR2X1 U57 ( .A(n17), .B(n87), .Y(n117) );
  XNOR2X1 U58 ( .A(n196), .B(n197), .Y(n108) );
  XOR2XL U59 ( .A(n18), .B(n192), .Y(n36) );
  XOR2XL U60 ( .A(n195), .B(n189), .Y(n58) );
  XNOR2X1 U61 ( .A(n17), .B(n197), .Y(n157) );
  XNOR2XL U62 ( .A(n142), .B(n83), .Y(P14[10]) );
  XOR2X1 U63 ( .A(n131), .B(n53), .Y(P9[4]) );
  XNOR2XL U64 ( .A(n94), .B(n86), .Y(n91) );
  XNOR2XL U65 ( .A(n20), .B(n117), .Y(P12[2]) );
  XOR2XL U66 ( .A(n107), .B(P1[2]), .Y(n55) );
  XNOR2XL U67 ( .A(n33), .B(n8), .Y(P6[10]) );
  XOR2XL U68 ( .A(n151), .B(n87), .Y(n52) );
  XOR2XL U69 ( .A(n123), .B(n124), .Y(P8[7]) );
  XNOR2XL U70 ( .A(P2[11]), .B(n5), .Y(P5[2]) );
  INVXL U71 ( .A(n188), .Y(n106) );
  INVXL U72 ( .A(n196), .Y(n20) );
  XNOR2XL U73 ( .A(n196), .B(n6), .Y(n45) );
  XNOR2XL U74 ( .A(n20), .B(n194), .Y(n40) );
  INVXL U75 ( .A(n191), .Y(n32) );
  XNOR2XL U76 ( .A(n17), .B(n189), .Y(n104) );
  XOR2X1 U77 ( .A(n14), .B(n134), .Y(n21) );
  XOR2X1 U78 ( .A(n195), .B(n191), .Y(n14) );
  XNOR2XL U79 ( .A(n199), .B(n193), .Y(n81) );
  XNOR2X1 U80 ( .A(n35), .B(n142), .Y(n92) );
  XNOR2XL U81 ( .A(n196), .B(n195), .Y(n35) );
  XNOR2XL U82 ( .A(n17), .B(n188), .Y(n76) );
  XOR2XL U83 ( .A(n196), .B(n188), .Y(n103) );
  XNOR2XL U84 ( .A(n18), .B(P1[2]), .Y(P12[12]) );
  XNOR2XL U85 ( .A(n120), .B(n6), .Y(P6[12]) );
  XNOR2X1 U86 ( .A(P5[2]), .B(n193), .Y(n65) );
  XNOR2XL U87 ( .A(P13[10]), .B(P1[12]), .Y(n115) );
  XOR2X1 U88 ( .A(n70), .B(n36), .Y(P4[10]) );
  XOR2X1 U89 ( .A(n131), .B(n44), .Y(n68) );
  XOR2XL U90 ( .A(n8), .B(n191), .Y(n44) );
  XOR2X1 U91 ( .A(n58), .B(n45), .Y(n98) );
  XNOR2XL U92 ( .A(n11), .B(n45), .Y(n88) );
  XNOR2XL U93 ( .A(n18), .B(n191), .Y(n141) );
  XNOR2XL U94 ( .A(n106), .B(n191), .Y(n133) );
  XOR2XL U95 ( .A(n4), .B(n154), .Y(n96) );
  XNOR2XL U96 ( .A(n195), .B(n6), .Y(n80) );
  XNOR2XL U97 ( .A(n18), .B(P12[11]), .Y(P2[12]) );
  XNOR2XL U98 ( .A(n187), .B(n90), .Y(P4[12]) );
  XOR2X1 U99 ( .A(n148), .B(n128), .Y(n137) );
  XNOR2XL U100 ( .A(n34), .B(n194), .Y(n148) );
  XNOR2XL U101 ( .A(n18), .B(n193), .Y(n102) );
  XNOR2XL U102 ( .A(n13), .B(P1[12]), .Y(P11[12]) );
  XNOR2XL U103 ( .A(n13), .B(n98), .Y(P2[6]) );
  XOR2X1 U104 ( .A(n110), .B(P6[2]), .Y(n101) );
  XOR2X1 U105 ( .A(n195), .B(b[9]), .Y(n110) );
  CLKBUFXL U106 ( .A(P12[5]), .Y(P13[0]) );
  XNOR2XL U107 ( .A(n199), .B(n109), .Y(P11[3]) );
  XNOR2XL U108 ( .A(n11), .B(n23), .Y(P9[3]) );
  XNOR2XL U109 ( .A(n190), .B(n74), .Y(P4[8]) );
  XNOR2XL U110 ( .A(n12), .B(n56), .Y(P6[6]) );
  CLKBUFXL U111 ( .A(P9[4]), .Y(P10[12]) );
  XNOR2XL U112 ( .A(P1[12]), .B(n126), .Y(P15[1]) );
  XNOR2X1 U113 ( .A(n20), .B(P12[12]), .Y(P2[0]) );
  XOR2X1 U114 ( .A(n145), .B(n28), .Y(P13[10]) );
  XNOR2X1 U115 ( .A(n13), .B(n129), .Y(P5[1]) );
  XNOR2X1 U116 ( .A(n42), .B(P1[1]), .Y(P12[11]) );
  XOR2X1 U117 ( .A(n122), .B(P6[10]), .Y(P16[0]) );
  XNOR2X1 U118 ( .A(n108), .B(n109), .Y(n23) );
  XNOR2X1 U119 ( .A(n63), .B(n74), .Y(P4[5]) );
  XNOR2X1 U120 ( .A(n122), .B(n137), .Y(P13[5]) );
  XNOR2X1 U121 ( .A(n136), .B(n137), .Y(P15[12]) );
  XNOR2X1 U122 ( .A(n5), .B(n69), .Y(P6[0]) );
  XNOR2X1 U123 ( .A(n12), .B(n112), .Y(P13[4]) );
  XOR2X1 U124 ( .A(n80), .B(n75), .Y(P5[12]) );
  XNOR2X1 U125 ( .A(n53), .B(n30), .Y(P11[2]) );
  XNOR2X1 U126 ( .A(n94), .B(n127), .Y(P1[3]) );
  XNOR2X1 U127 ( .A(n8), .B(n122), .Y(n154) );
  XNOR2X1 U128 ( .A(n199), .B(n66), .Y(n27) );
  XNOR2X1 U129 ( .A(n9), .B(n76), .Y(n143) );
  XNOR2X1 U130 ( .A(n54), .B(n134), .Y(n105) );
  XNOR2X1 U131 ( .A(n199), .B(P1[2]), .Y(n129) );
  XNOR2X1 U132 ( .A(n48), .B(n12), .Y(n60) );
  XOR2X1 U133 ( .A(n23), .B(n107), .Y(P8[2]) );
  XOR2X1 U134 ( .A(n116), .B(n134), .Y(n84) );
  XOR2X1 U135 ( .A(n116), .B(n118), .Y(n69) );
  XOR2X1 U136 ( .A(n147), .B(P1[11]), .Y(n124) );
  XOR2X1 U137 ( .A(n89), .B(n13), .Y(P13[8]) );
  XOR2X1 U138 ( .A(n103), .B(n124), .Y(n86) );
  XOR2X1 U139 ( .A(n90), .B(n8), .Y(P13[7]) );
  XOR2X1 U140 ( .A(n78), .B(n79), .Y(n74) );
  XNOR2X1 U141 ( .A(n53), .B(P8[2]), .Y(P16[6]) );
  XNOR2X1 U142 ( .A(n106), .B(P13[7]), .Y(P16[7]) );
  XNOR2X1 U143 ( .A(n61), .B(P13[8]), .Y(P16[8]) );
  XNOR2X1 U144 ( .A(n10), .B(n111), .Y(P16[4]) );
  XNOR2X1 U145 ( .A(n6), .B(P4[10]), .Y(P16[5]) );
  XNOR2X1 U146 ( .A(P12[5]), .B(n116), .Y(n78) );
  XNOR2XL U147 ( .A(n145), .B(n42), .Y(n89) );
  XNOR2X1 U148 ( .A(P1[7]), .B(n129), .Y(n90) );
  XOR2X1 U149 ( .A(n87), .B(n41), .Y(P3[6]) );
  XNOR2X1 U150 ( .A(n56), .B(n30), .Y(n48) );
  XOR2X1 U151 ( .A(P9[0]), .B(n146), .Y(n112) );
  XNOR2X1 U152 ( .A(n135), .B(n143), .Y(n29) );
  XOR2X1 U153 ( .A(P11[7]), .B(n66), .Y(n59) );
  XOR2X1 U154 ( .A(n138), .B(n152), .Y(n139) );
  XNOR2X1 U155 ( .A(n199), .B(n104), .Y(n152) );
  XNOR2X1 U156 ( .A(P9[4]), .B(n8), .Y(P4[1]) );
  XNOR2X1 U157 ( .A(n6), .B(n160), .Y(P10[5]) );
  XNOR2X1 U158 ( .A(n5), .B(n147), .Y(P6[2]) );
  XOR2X1 U159 ( .A(n127), .B(P11[11]), .Y(n22) );
  XOR2X1 U160 ( .A(n63), .B(P8[7]), .Y(P16[12]) );
  XNOR2X1 U161 ( .A(n1), .B(n40), .Y(P11[5]) );
  XNOR2X1 U162 ( .A(n5), .B(n21), .Y(P9[12]) );
  XNOR2X1 U163 ( .A(n13), .B(n43), .Y(P8[0]) );
  XNOR2X1 U164 ( .A(n10), .B(n59), .Y(P7[12]) );
  XNOR2X1 U165 ( .A(n8), .B(n99), .Y(P3[0]) );
  XNOR2X1 U166 ( .A(n10), .B(n100), .Y(P3[12]) );
  XOR2X1 U167 ( .A(P11[11]), .B(n57), .Y(P7[0]) );
  XNOR2X1 U168 ( .A(n1), .B(n63), .Y(n31) );
  XNOR2X1 U169 ( .A(n61), .B(n92), .Y(n85) );
  XNOR2X1 U170 ( .A(n10), .B(n95), .Y(P6[1]) );
  XNOR2X1 U171 ( .A(n108), .B(P10[5]), .Y(n19) );
  XOR2X1 U172 ( .A(P11[11]), .B(n52), .Y(n121) );
  XOR2X1 U173 ( .A(P1[1]), .B(n45), .Y(P6[8]) );
  XOR2X1 U174 ( .A(n46), .B(n47), .Y(n43) );
  XNOR2X1 U175 ( .A(n53), .B(n63), .Y(n99) );
  XNOR2X1 U176 ( .A(n94), .B(n107), .Y(n151) );
  XNOR2X1 U177 ( .A(n199), .B(n97), .Y(n39) );
  XNOR2X1 U178 ( .A(n10), .B(n92), .Y(n113) );
  XNOR2X1 U179 ( .A(n17), .B(P6[8]), .Y(n16) );
  XNOR2X1 U180 ( .A(n18), .B(n190), .Y(n134) );
  XNOR2X1 U181 ( .A(n197), .B(n42), .Y(n87) );
  XOR2X1 U182 ( .A(n196), .B(n51), .Y(P11[7]) );
  XNOR2X1 U183 ( .A(P9[5]), .B(n190), .Y(n83) );
  XOR2X1 U184 ( .A(n195), .B(n29), .Y(P9[5]) );
  XNOR2X1 U185 ( .A(n17), .B(n190), .Y(P1[11]) );
  XNOR2X1 U186 ( .A(n192), .B(n9), .Y(P1[1]) );
  XNOR2X1 U187 ( .A(n188), .B(n61), .Y(n66) );
  XOR2X1 U188 ( .A(n194), .B(P11[7]), .Y(P2[2]) );
  XOR2X1 U189 ( .A(n196), .B(n191), .Y(n122) );
  XNOR2X1 U190 ( .A(n130), .B(n83), .Y(P15[0]) );
  XNOR2X1 U191 ( .A(n188), .B(n48), .Y(P8[12]) );
  XNOR2X1 U192 ( .A(n188), .B(n89), .Y(P4[0]) );
  XNOR2X1 U193 ( .A(n53), .B(n191), .Y(n79) );
  XNOR2X1 U194 ( .A(n11), .B(n87), .Y(P11[6]) );
  XNOR2X1 U195 ( .A(n111), .B(n4), .Y(n73) );
  XOR2X1 U196 ( .A(n130), .B(n160), .Y(n150) );
  XOR2X1 U197 ( .A(P3[7]), .B(n81), .Y(n75) );
  XOR2X1 U198 ( .A(P3[6]), .B(n77), .Y(n71) );
  XNOR2X1 U199 ( .A(n197), .B(n72), .Y(P16[3]) );
  XNOR2X1 U200 ( .A(n190), .B(n115), .Y(P16[1]) );
  XNOR2X1 U201 ( .A(n188), .B(n115), .Y(P16[10]) );
  XNOR2X1 U202 ( .A(b[6]), .B(n105), .Y(P16[9]) );
  XNOR2X1 U203 ( .A(n197), .B(n53), .Y(n147) );
  XNOR2X1 U204 ( .A(n194), .B(n42), .Y(n127) );
  XNOR2X1 U205 ( .A(n25), .B(n141), .Y(n38) );
  XOR2X1 U206 ( .A(n195), .B(n84), .Y(P7[2]) );
  XOR2X1 U207 ( .A(n187), .B(n134), .Y(n138) );
  XNOR2X1 U208 ( .A(n125), .B(n187), .Y(n25) );
  XNOR2X1 U209 ( .A(n197), .B(n32), .Y(n142) );
  XNOR2X1 U210 ( .A(P10[2]), .B(n4), .Y(n50) );
  XNOR2X1 U211 ( .A(P2[10]), .B(P1[0]), .Y(n67) );
  XOR2X1 U212 ( .A(n4), .B(P11[6]), .Y(P1[7]) );
  XOR2X1 U213 ( .A(n191), .B(P1[3]), .Y(P2[11]) );
  XOR2X1 U214 ( .A(n194), .B(n154), .Y(P10[2]) );
  XOR2X1 U215 ( .A(n4), .B(P5[1]), .Y(P2[10]) );
  XOR2X1 U216 ( .A(n194), .B(n100), .Y(n33) );
  XOR2X1 U217 ( .A(n187), .B(n92), .Y(n54) );
  XOR2X1 U218 ( .A(n191), .B(n117), .Y(n56) );
  XOR2X1 U219 ( .A(n4), .B(P11[2]), .Y(n125) );
  XOR2X1 U220 ( .A(P7[2]), .B(n133), .Y(n111) );
  INVX1 U221 ( .A(n197), .Y(n28) );
  XNOR2X1 U222 ( .A(n194), .B(n189), .Y(n135) );
  XOR2X1 U223 ( .A(n192), .B(n79), .Y(P12[10]) );
  XOR2X1 U224 ( .A(n47), .B(n88), .Y(n41) );
  INVX1 U225 ( .A(n189), .Y(n61) );
  XNOR2X1 U226 ( .A(P2[2]), .B(n192), .Y(n145) );
  BUFX3 U227 ( .A(n32), .Y(n199) );
  XNOR2X1 U228 ( .A(n188), .B(n18), .Y(n63) );
  XNOR2X1 U229 ( .A(n189), .B(n12), .Y(P11[11]) );
  XNOR2X1 U230 ( .A(n187), .B(n106), .Y(n107) );
  XOR2X1 U231 ( .A(n99), .B(n157), .Y(P13[12]) );
  XNOR2X1 U232 ( .A(n93), .B(n31), .Y(n62) );
  XNOR2X1 U233 ( .A(n187), .B(n190), .Y(n93) );
  XNOR2X1 U234 ( .A(n187), .B(n18), .Y(n128) );
  XNOR2X1 U235 ( .A(n96), .B(n192), .Y(n82) );
  XOR2X1 U236 ( .A(n113), .B(n114), .Y(P16[2]) );
  XNOR2X1 U237 ( .A(n17), .B(n192), .Y(n114) );
  XNOR2X1 U238 ( .A(n1), .B(n190), .Y(n140) );
  XNOR2X1 U239 ( .A(n42), .B(n193), .Y(n146) );
  XNOR2X1 U240 ( .A(n20), .B(n4), .Y(n95) );
  XOR2X1 U241 ( .A(n192), .B(n51), .Y(n46) );
  XNOR2X1 U242 ( .A(n195), .B(n106), .Y(n136) );
  XNOR2X1 U243 ( .A(n196), .B(n190), .Y(n24) );
  XOR2X1 U244 ( .A(n196), .B(b[9]), .Y(n130) );
  XNOR2X1 U245 ( .A(n7), .B(n71), .Y(P5[11]) );
  XNOR2X1 U246 ( .A(P6[12]), .B(n119), .Y(P15[7]) );
  XNOR2X1 U247 ( .A(n7), .B(n138), .Y(P14[3]) );
  XOR2X1 U248 ( .A(b[9]), .B(n86), .Y(P3[7]) );
  XOR2X1 U249 ( .A(b[9]), .B(n118), .Y(n120) );
  BUFX3 U250 ( .A(b[4]), .Y(n191) );
  XNOR2X1 U251 ( .A(n53), .B(n69), .Y(P15[8]) );
  XOR2X1 U252 ( .A(n135), .B(n105), .Y(P14[6]) );
  XNOR2X1 U253 ( .A(n11), .B(n57), .Y(P12[1]) );
  XOR2X1 U254 ( .A(n95), .B(n101), .Y(P12[3]) );
  XNOR2X1 U255 ( .A(n106), .B(n81), .Y(P11[1]) );
  XOR2X1 U256 ( .A(n134), .B(n143), .Y(P10[1]) );
  XNOR2X1 U258 ( .A(n8), .B(n55), .Y(P10[7]) );
  XNOR2X1 U259 ( .A(n106), .B(n22), .Y(P10[8]) );
  XOR2X1 U260 ( .A(n26), .B(n27), .Y(P9[1]) );
  XNOR2X1 U261 ( .A(n20), .B(n21), .Y(P9[7]) );
  XNOR2X1 U262 ( .A(n20), .B(n38), .Y(P8[1]) );
  XNOR2X1 U263 ( .A(n8), .B(n62), .Y(P6[11]) );
  XOR2X1 U264 ( .A(n76), .B(n71), .Y(P4[6]) );
  XNOR2X1 U265 ( .A(n7), .B(n23), .Y(P4[11]) );
  XNOR2X1 U266 ( .A(n94), .B(P6[2]), .Y(P3[11]) );
  XNOR2X1 U267 ( .A(n11), .B(n39), .Y(P2[7]) );
  XNOR2X1 U268 ( .A(n94), .B(n120), .Y(P14[2]) );
  XNOR2X1 U269 ( .A(n106), .B(n125), .Y(P15[2]) );
  XNOR2X1 U270 ( .A(n20), .B(n49), .Y(P13[2]) );
  XNOR2X1 U271 ( .A(n199), .B(n121), .Y(P13[3]) );
  XOR2X1 U272 ( .A(n146), .B(n91), .Y(P13[6]) );
  XOR2X1 U273 ( .A(n123), .B(P12[2]), .Y(P13[11]) );
  XOR2X1 U274 ( .A(n51), .B(n52), .Y(P7[11]) );
  XNOR2X1 U275 ( .A(n7), .B(n54), .Y(P7[10]) );
  XNOR2X1 U276 ( .A(n45), .B(n73), .Y(P14[7]) );
  XNOR2X1 U277 ( .A(n67), .B(n128), .Y(P15[10]) );
  XNOR2X1 U278 ( .A(n106), .B(n96), .Y(P12[7]) );
  XNOR2X1 U279 ( .A(n11), .B(n121), .Y(P15[6]) );
  XNOR2X1 U280 ( .A(n1), .B(n43), .Y(P7[8]) );
  XNOR2X1 U281 ( .A(n199), .B(n33), .Y(P8[8]) );
  XNOR2X1 U282 ( .A(n199), .B(n46), .Y(P6[7]) );
  XOR2X1 U283 ( .A(n130), .B(n68), .Y(P14[8]) );
  XNOR2X1 U284 ( .A(n11), .B(n19), .Y(P9[8]) );
  XNOR2X1 U285 ( .A(n106), .B(n104), .Y(P11[10]) );
  XOR2X1 U286 ( .A(n38), .B(n140), .Y(P14[11]) );
  XNOR2X1 U287 ( .A(n11), .B(n97), .Y(P12[6]) );
  XNOR2X1 U288 ( .A(n20), .B(n34), .Y(P8[6]) );
  XNOR2X1 U289 ( .A(n13), .B(n149), .Y(P12[8]) );
  XNOR2X1 U290 ( .A(n11), .B(n22), .Y(P9[6]) );
  XNOR2X1 U291 ( .A(n10), .B(n19), .Y(P10[11]) );
  XOR2X1 U292 ( .A(P1[11]), .B(n81), .Y(P12[9]) );
  XNOR2X1 U293 ( .A(n10), .B(n151), .Y(P10[6]) );
  XNOR2X1 U294 ( .A(n66), .B(n67), .Y(P5[7]) );
  XNOR2X1 U295 ( .A(n12), .B(n68), .Y(P5[6]) );
  XNOR2X1 U296 ( .A(n65), .B(n103), .Y(P15[11]) );
  XNOR2X1 U297 ( .A(n11), .B(n113), .Y(P13[9]) );
  XOR2X1 U298 ( .A(n39), .B(n40), .Y(P8[11]) );
  XNOR2X1 U299 ( .A(n196), .B(n60), .Y(P6[3]) );
  XNOR2X1 U300 ( .A(n12), .B(P2[0]), .Y(P7[9]) );
  XNOR2X1 U301 ( .A(n1), .B(n37), .Y(P7[7]) );
  XNOR2X1 U302 ( .A(n13), .B(n37), .Y(P8[3]) );
  XNOR2X1 U303 ( .A(n8), .B(n75), .Y(P4[7]) );
  XOR2X1 U304 ( .A(n24), .B(n25), .Y(P9[2]) );
  XNOR2X1 U305 ( .A(n106), .B(P2[2]), .Y(P15[3]) );
  XNOR2X1 U306 ( .A(n189), .B(n64), .Y(P5[8]) );
  XNOR2X1 U307 ( .A(n63), .B(n64), .Y(P5[9]) );
  XNOR2X1 U308 ( .A(n8), .B(n21), .Y(P10[9]) );
  XNOR2X1 U309 ( .A(n194), .B(n72), .Y(P5[10]) );
  XNOR2X1 U310 ( .A(n187), .B(n83), .Y(P4[2]) );
  XNOR2X1 U311 ( .A(n12), .B(n150), .Y(P10[10]) );
  XNOR2X1 U312 ( .A(n195), .B(n50), .Y(P7[1]) );
  XOR2X1 U313 ( .A(P1[2]), .B(n49), .Y(P7[3]) );
  XNOR2X1 U314 ( .A(n197), .B(n70), .Y(P5[3]) );
  XOR2X1 U315 ( .A(n63), .B(n85), .Y(P3[2]) );
  XNOR2X1 U316 ( .A(n5), .B(n91), .Y(P3[3]) );
  XNOR2X1 U317 ( .A(n17), .B(n85), .Y(P3[8]) );
  XNOR2X1 U318 ( .A(n17), .B(n84), .Y(P3[9]) );
  XNOR2X1 U319 ( .A(n199), .B(P6[1]), .Y(P3[10]) );
  XNOR2X1 U320 ( .A(n1), .B(n26), .Y(P2[1]) );
  XNOR2X1 U321 ( .A(n10), .B(n101), .Y(P2[3]) );
  XNOR2X1 U322 ( .A(n188), .B(n82), .Y(P2[8]) );
  XNOR2X1 U323 ( .A(n5), .B(P11[7]), .Y(P1[8]) );
  XOR2X1 U324 ( .A(n139), .B(n136), .Y(P14[1]) );
  XOR2X1 U325 ( .A(n140), .B(n153), .Y(P13[1]) );
  INVX1 U326 ( .A(b[9]), .Y(n18) );
  BUFX3 U327 ( .A(b[6]), .Y(n193) );
  BUFX3 U328 ( .A(b_3), .Y(n190) );
  BUFX3 U329 ( .A(b_2), .Y(n189) );
  BUFX3 U330 ( .A(b[7]), .Y(n194) );
  XNOR2X1 U331 ( .A(b[6]), .B(n60), .Y(P15[9]) );
  XNOR2X1 U332 ( .A(n190), .B(n82), .Y(P4[3]) );
  XNOR2X1 U333 ( .A(b[6]), .B(n73), .Y(P4[9]) );
  XOR2X1 U334 ( .A(n30), .B(n31), .Y(P8[9]) );
  XOR2X1 U335 ( .A(n40), .B(n62), .Y(P3[1]) );
  BUFX3 U336 ( .A(P9[0]), .Y(P8[5]) );
  BUFX3 U337 ( .A(P16[12]), .Y(P15[4]) );
  BUFX3 U338 ( .A(P9[5]), .Y(P10[0]) );
  BUFX3 U339 ( .A(P6[12]), .Y(P5[4]) );
  BUFX3 U340 ( .A(P13[12]), .Y(P12[4]) );
  BUFX3 U341 ( .A(P8[12]), .Y(P7[4]) );
  BUFX3 U342 ( .A(P4[5]), .Y(P5[0]) );
  BUFX3 U343 ( .A(P6[0]), .Y(P5[5]) );
  BUFX3 U344 ( .A(P4[0]), .Y(P3[5]) );
  BUFX3 U345 ( .A(P3[12]), .Y(P2[4]) );
  BUFX3 U346 ( .A(P15[0]), .Y(P14[5]) );
  BUFX3 U347 ( .A(P7[12]), .Y(P6[4]) );
  BUFX3 U348 ( .A(P9[12]), .Y(P8[4]) );
  BUFX3 U349 ( .A(P13[4]), .Y(P14[12]) );
  BUFX3 U350 ( .A(P7[0]), .Y(P6[5]) );
  BUFX3 U351 ( .A(P4[12]), .Y(P3[4]) );
  BUFX3 U352 ( .A(P11[12]), .Y(P10[4]) );
  BUFX3 U353 ( .A(P15[12]), .Y(P14[4]) );
  BUFX3 U354 ( .A(P8[0]), .Y(P7[5]) );
  BUFX3 U355 ( .A(P3[0]), .Y(P2[5]) );
  BUFX3 U356 ( .A(P2[12]), .Y(P1[4]) );
  BUFX3 U357 ( .A(b[10]), .Y(n196) );
  BUFX3 U358 ( .A(P11[5]), .Y(P12[0]) );
  BUFX3 U359 ( .A(P12[12]), .Y(P11[4]) );
  BUFX3 U360 ( .A(P13[5]), .Y(P14[0]) );
  BUFX3 U361 ( .A(P10[5]), .Y(P11[0]) );
  BUFX3 U362 ( .A(P2[0]), .Y(P1[5]) );
  BUFX3 U363 ( .A(P5[12]), .Y(P4[4]) );
  XOR2X1 U364 ( .A(n15), .B(n16), .Y(P9[9]) );
  XNOR2X1 U365 ( .A(n28), .B(n29), .Y(P9[10]) );
  XNOR2X1 U366 ( .A(n132), .B(n55), .Y(P6[9]) );
  XNOR2X1 U367 ( .A(n28), .B(n103), .Y(P1[9]) );
  XNOR2X1 U368 ( .A(n28), .B(P11[5]), .Y(P1[6]) );
  XNOR2X1 U369 ( .A(n132), .B(n104), .Y(P1[10]) );
  XNOR2X1 U370 ( .A(n28), .B(n59), .Y(n153) );
  XOR2XL U371 ( .A(P12[10]), .B(n15), .Y(n37) );
  XNOR2X1 U372 ( .A(n28), .B(n102), .Y(n26) );
  XNOR2X1 U373 ( .A(n28), .B(n139), .Y(n49) );
  XNOR2X1 U374 ( .A(n28), .B(n40), .Y(n57) );
  XNOR2X1 U375 ( .A(n28), .B(n30), .Y(n149) );
endmodule


module multiplier_column7_p16 ( b, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, 
        P11, P12, P13, P14, P15, P16 );
  input [12:0] b;
  output [12:0] P1;
  output [12:0] P2;
  output [12:0] P3;
  output [12:0] P4;
  output [12:0] P5;
  output [12:0] P6;
  output [12:0] P7;
  output [12:0] P8;
  output [12:0] P9;
  output [12:0] P10;
  output [12:0] P11;
  output [12:0] P12;
  output [12:0] P13;
  output [12:0] P14;
  output [12:0] P15;
  output [12:0] P16;
  wire   b_3, b_2, b_1, b_0, n210, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n76, n77, n78, n79, n80, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n132, n133, n134, n136, n137,
         n138, n139, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n32, n47, n61, n75, n81, n103,
         n131, n135, n140, n156, n157, n158, n159, n207;
  assign b_3 = b[3];
  assign b_2 = b[2];
  assign b_1 = b[1];
  assign b_0 = b[0];

  XNOR2X4 U279 ( .A(b[4]), .B(n23), .Y(n77) );
  XOR2X1 U1 ( .A(b[9]), .B(P13[12]), .Y(P2[2]) );
  XNOR2X2 U2 ( .A(P7[4]), .B(n86), .Y(n80) );
  XNOR2XL U3 ( .A(n49), .B(n50), .Y(P8[4]) );
  XNOR2X2 U4 ( .A(n21), .B(n50), .Y(n110) );
  XNOR2X2 U5 ( .A(n102), .B(n77), .Y(n57) );
  XNOR2X2 U6 ( .A(n45), .B(n210), .Y(P13[8]) );
  XNOR2X2 U7 ( .A(n54), .B(b[8]), .Y(n210) );
  BUFX3 U8 ( .A(P15[6]), .Y(P16[0]) );
  CLKINVXL U9 ( .A(b[10]), .Y(n13) );
  INVX2 U10 ( .A(b[11]), .Y(n113) );
  CLKINVXL U11 ( .A(b[11]), .Y(n135) );
  XNOR2X2 U12 ( .A(n118), .B(n125), .Y(n33) );
  INVX8 U13 ( .A(b[10]), .Y(n45) );
  XNOR2X4 U14 ( .A(b[8]), .B(n48), .Y(n137) );
  INVX4 U15 ( .A(b[9]), .Y(n48) );
  INVX1 U16 ( .A(n77), .Y(n150) );
  XNOR2X1 U17 ( .A(P12[4]), .B(n150), .Y(n149) );
  CLKBUFX8 U18 ( .A(b[12]), .Y(n207) );
  BUFX3 U19 ( .A(n105), .Y(n1) );
  INVX1 U20 ( .A(n76), .Y(n144) );
  XNOR2X1 U21 ( .A(n119), .B(n133), .Y(n124) );
  XOR2X1 U22 ( .A(P1[0]), .B(n149), .Y(P11[8]) );
  XOR2X1 U23 ( .A(P2[2]), .B(n90), .Y(P7[4]) );
  XNOR2X1 U24 ( .A(n39), .B(n137), .Y(P1[3]) );
  XOR2X1 U25 ( .A(b[5]), .B(P1[3]), .Y(P2[10]) );
  XOR2X1 U26 ( .A(n33), .B(n44), .Y(n66) );
  XOR2X1 U27 ( .A(P1[11]), .B(n110), .Y(n117) );
  XNOR2X1 U28 ( .A(n22), .B(n124), .Y(P16[9]) );
  XOR2X1 U29 ( .A(P11[8]), .B(n4), .Y(n111) );
  OAI2BB1X2 U30 ( .A0N(n15), .A1N(n51), .B0(n16), .Y(n108) );
  INVX1 U31 ( .A(P8[10]), .Y(n15) );
  XOR2X1 U32 ( .A(n76), .B(n105), .Y(P13[12]) );
  XOR2X1 U33 ( .A(n137), .B(P1[8]), .Y(n123) );
  OAI2BB1X1 U34 ( .A0N(n136), .A1N(n54), .B0(n61), .Y(P12[3]) );
  XNOR2XL U35 ( .A(b_0), .B(n3), .Y(n22) );
  XNOR2X2 U36 ( .A(b_0), .B(n30), .Y(n76) );
  XNOR2XL U37 ( .A(n3), .B(b[10]), .Y(n62) );
  XNOR2X1 U38 ( .A(b[10]), .B(b_1), .Y(n145) );
  XOR2XL U39 ( .A(P1[0]), .B(b[10]), .Y(n159) );
  XOR2XL U40 ( .A(n54), .B(b[10]), .Y(n158) );
  XNOR2X4 U41 ( .A(b[11]), .B(n45), .Y(n29) );
  XOR2X2 U42 ( .A(n43), .B(n64), .Y(n87) );
  XNOR2X1 U43 ( .A(P2[10]), .B(b_2), .Y(n43) );
  CLKINVX3 U44 ( .A(b[5]), .Y(n23) );
  XNOR2X1 U45 ( .A(b[11]), .B(n14), .Y(n105) );
  INVX1 U46 ( .A(b[12]), .Y(n14) );
  XNOR2X1 U47 ( .A(b_2), .B(n48), .Y(n114) );
  XOR2X1 U48 ( .A(n109), .B(n1), .Y(n132) );
  XOR2X2 U49 ( .A(b_0), .B(n29), .Y(P12[4]) );
  XNOR2X1 U50 ( .A(n114), .B(n111), .Y(P15[6]) );
  CLKINVX3 U51 ( .A(b[7]), .Y(n54) );
  INVX1 U52 ( .A(b[7]), .Y(n4) );
  XNOR2X2 U53 ( .A(P1[0]), .B(n102), .Y(n96) );
  INVX4 U54 ( .A(n207), .Y(n102) );
  XNOR2XL U55 ( .A(n54), .B(n55), .Y(P8[1]) );
  XNOR2X1 U56 ( .A(P14[11]), .B(n54), .Y(P2[8]) );
  BUFX3 U57 ( .A(P14[11]), .Y(P13[4]) );
  XOR2X2 U58 ( .A(n207), .B(n91), .Y(P14[11]) );
  XNOR2XL U59 ( .A(n6), .B(n27), .Y(P7[10]) );
  XNOR2X4 U60 ( .A(n113), .B(b_1), .Y(n44) );
  XNOR2X1 U61 ( .A(b_3), .B(P1[8]), .Y(n68) );
  XNOR2XL U62 ( .A(n207), .B(n43), .Y(P8[8]) );
  XNOR2X1 U63 ( .A(n135), .B(n92), .Y(n64) );
  INVX1 U64 ( .A(b_0), .Y(n70) );
  INVX1 U65 ( .A(b_3), .Y(n42) );
  INVX4 U66 ( .A(b_1), .Y(n30) );
  CLKINVX3 U67 ( .A(n83), .Y(n21) );
  XOR2X1 U68 ( .A(n156), .B(n132), .Y(n100) );
  XNOR2X1 U69 ( .A(P12[0]), .B(n207), .Y(n95) );
  XNOR2X1 U70 ( .A(n84), .B(n85), .Y(n82) );
  BUFX3 U71 ( .A(n48), .Y(n12) );
  INVX1 U72 ( .A(n210), .Y(n17) );
  BUFX3 U73 ( .A(n30), .Y(n6) );
  XNOR2X1 U74 ( .A(n10), .B(n100), .Y(n52) );
  INVX1 U75 ( .A(b_0), .Y(n10) );
  INVX1 U76 ( .A(b_3), .Y(n7) );
  BUFX8 U77 ( .A(b[6]), .Y(P1[0]) );
  INVX1 U78 ( .A(b[4]), .Y(n25) );
  INVX1 U79 ( .A(b[5]), .Y(n11) );
  BUFX3 U80 ( .A(P6[0]), .Y(P5[6]) );
  XNOR2X1 U81 ( .A(n3), .B(n100), .Y(n34) );
  XNOR2X1 U82 ( .A(n51), .B(P1[2]), .Y(n152) );
  INVX1 U83 ( .A(n4), .Y(n5) );
  XOR2X1 U84 ( .A(n65), .B(n127), .Y(P16[10]) );
  XOR2X1 U85 ( .A(P1[5]), .B(n69), .Y(P8[10]) );
  BUFX3 U86 ( .A(P1[5]), .Y(P2[12]) );
  XOR2X2 U87 ( .A(b[11]), .B(P13[8]), .Y(P1[5]) );
  XNOR2X1 U88 ( .A(n107), .B(n108), .Y(P4[4]) );
  XNOR2X2 U89 ( .A(n45), .B(n44), .Y(P1[8]) );
  XOR2X1 U90 ( .A(P2[8]), .B(n128), .Y(n65) );
  XOR2X4 U91 ( .A(n106), .B(n13), .Y(P16[12]) );
  XNOR2X2 U92 ( .A(n117), .B(n142), .Y(n106) );
  XNOR2X1 U93 ( .A(n10), .B(P16[12]), .Y(P11[3]) );
  XNOR2X1 U94 ( .A(b[7]), .B(n48), .Y(n109) );
  XOR2X1 U95 ( .A(P1[11]), .B(P13[0]), .Y(n121) );
  XNOR2X2 U96 ( .A(n86), .B(n87), .Y(P6[0]) );
  XNOR2XL U97 ( .A(n13), .B(P1[3]), .Y(P14[2]) );
  CLKBUFX2 U98 ( .A(b[4]), .Y(P1[11]) );
  XNOR2X2 U99 ( .A(b[4]), .B(n21), .Y(n91) );
  INVX1 U100 ( .A(b_2), .Y(n3) );
  XNOR2XL U101 ( .A(n3), .B(n84), .Y(P15[1]) );
  XNOR2XL U102 ( .A(n3), .B(n123), .Y(P2[3]) );
  XNOR2XL U103 ( .A(n3), .B(n1), .Y(P1[9]) );
  INVX1 U104 ( .A(b_2), .Y(n74) );
  XNOR2X1 U105 ( .A(b_2), .B(n30), .Y(n128) );
  XNOR2XL U106 ( .A(n7), .B(b_0), .Y(n72) );
  INVX1 U107 ( .A(b[8]), .Y(n9) );
  INVX1 U108 ( .A(b[8]), .Y(n8) );
  XNOR2XL U109 ( .A(n8), .B(n76), .Y(n40) );
  XNOR2XL U110 ( .A(n10), .B(n77), .Y(P12[9]) );
  XNOR2XL U111 ( .A(n10), .B(n97), .Y(P15[3]) );
  XNOR2XL U112 ( .A(n121), .B(n11), .Y(P6[1]) );
  XNOR2XL U113 ( .A(n11), .B(n5), .Y(n133) );
  XNOR2X1 U114 ( .A(n23), .B(b[9]), .Y(n142) );
  XNOR2XL U115 ( .A(n45), .B(b[9]), .Y(n19) );
  XNOR2X1 U116 ( .A(n102), .B(n128), .Y(P13[0]) );
  XNOR2XL U117 ( .A(n9), .B(b[11]), .Y(n127) );
  XNOR2X1 U118 ( .A(n39), .B(P12[3]), .Y(P16[5]) );
  XNOR2X1 U119 ( .A(n144), .B(P1[10]), .Y(n143) );
  XNOR2X1 U120 ( .A(n6), .B(P1[10]), .Y(P13[1]) );
  NAND2X1 U121 ( .A(P8[10]), .B(P12[7]), .Y(n16) );
  INVX1 U122 ( .A(n17), .Y(P1[2]) );
  NAND2X1 U123 ( .A(n32), .B(n47), .Y(n61) );
  INVX1 U124 ( .A(n136), .Y(n32) );
  INVXL U125 ( .A(n54), .Y(n47) );
  XNOR2X1 U126 ( .A(n145), .B(n146), .Y(n136) );
  CLKBUFX2 U127 ( .A(P3[4]), .Y(P4[11]) );
  XOR2X1 U128 ( .A(P12[8]), .B(n137), .Y(n151) );
  XOR2X1 U129 ( .A(n92), .B(n123), .Y(n84) );
  XNOR2X1 U130 ( .A(n6), .B(n132), .Y(P15[0]) );
  XNOR2X1 U131 ( .A(b[8]), .B(n124), .Y(P15[7]) );
  XOR2XL U132 ( .A(n109), .B(n110), .Y(P4[3]) );
  XNOR2X1 U133 ( .A(n25), .B(n26), .Y(P9[7]) );
  BUFX2 U134 ( .A(P3[6]), .Y(P4[0]) );
  BUFX2 U135 ( .A(P2[0]), .Y(P1[6]) );
  XOR2X1 U136 ( .A(n91), .B(n92), .Y(n46) );
  XOR2X1 U137 ( .A(n97), .B(n98), .Y(P7[3]) );
  XOR2X1 U138 ( .A(n19), .B(n66), .Y(P16[8]) );
  CLKBUFXL U139 ( .A(P15[0]), .Y(P14[6]) );
  CLKBUFXL U140 ( .A(P16[12]), .Y(P15[5]) );
  XNOR2X1 U141 ( .A(n68), .B(n96), .Y(n119) );
  XNOR2X1 U142 ( .A(n8), .B(P12[4]), .Y(P2[1]) );
  XNOR2XL U143 ( .A(n39), .B(n47), .Y(P1[1]) );
  XNOR2XL U144 ( .A(n10), .B(n102), .Y(n94) );
  INVX8 U145 ( .A(P1[0]), .Y(n39) );
  XNOR2X1 U146 ( .A(n113), .B(b[9]), .Y(n98) );
  XNOR2XL U147 ( .A(P2[1]), .B(n114), .Y(n78) );
  XNOR2XL U148 ( .A(n30), .B(n73), .Y(n24) );
  XNOR2X1 U149 ( .A(P13[2]), .B(n75), .Y(n126) );
  XOR2X1 U150 ( .A(n30), .B(n86), .Y(n75) );
  XNOR2X1 U151 ( .A(n11), .B(n65), .Y(P6[9]) );
  XNOR2X1 U152 ( .A(b[8]), .B(n30), .Y(n50) );
  XNOR2X1 U153 ( .A(n8), .B(n34), .Y(P15[8]) );
  XNOR2XL U154 ( .A(n135), .B(P1[11]), .Y(n138) );
  CLKBUFXL U155 ( .A(P13[12]), .Y(P12[5]) );
  CLKBUFXL U156 ( .A(P12[0]), .Y(P11[6]) );
  XOR2X1 U157 ( .A(n5), .B(n126), .Y(n97) );
  XNOR2XL U158 ( .A(n12), .B(n57), .Y(P7[8]) );
  XNOR2XL U159 ( .A(n10), .B(n151), .Y(P10[10]) );
  XOR2X1 U160 ( .A(n72), .B(n122), .Y(P2[4]) );
  XOR2X1 U161 ( .A(n79), .B(n89), .Y(P5[4]) );
  XOR2X1 U162 ( .A(P10[2]), .B(n134), .Y(P15[4]) );
  XOR2X1 U163 ( .A(n81), .B(n107), .Y(n99) );
  XNOR2XL U164 ( .A(b_1), .B(P13[8]), .Y(n81) );
  XOR2X1 U165 ( .A(n132), .B(n103), .Y(P15[11]) );
  XNOR2XL U166 ( .A(n13), .B(b[5]), .Y(n103) );
  XNOR2X1 U167 ( .A(n80), .B(n131), .Y(P5[9]) );
  XOR2X1 U168 ( .A(P1[0]), .B(b_2), .Y(n131) );
  XOR2X1 U169 ( .A(n159), .B(n104), .Y(n88) );
  CLKBUFXL U170 ( .A(b[5]), .Y(P1[12]) );
  BUFX3 U171 ( .A(P11[0]), .Y(P10[6]) );
  BUFX3 U172 ( .A(P4[5]), .Y(P5[12]) );
  BUFX3 U173 ( .A(P10[0]), .Y(P9[6]) );
  BUFX3 U174 ( .A(P11[11]), .Y(P10[4]) );
  BUFX3 U175 ( .A(P15[12]), .Y(P14[5]) );
  XNOR2X1 U176 ( .A(n150), .B(n19), .Y(n31) );
  XOR2XL U177 ( .A(n28), .B(n29), .Y(P10[12]) );
  XOR2X1 U178 ( .A(P1[10]), .B(n27), .Y(P10[0]) );
  XNOR2X1 U179 ( .A(n135), .B(n55), .Y(P4[12]) );
  XNOR2X1 U180 ( .A(n12), .B(n152), .Y(P11[11]) );
  XNOR2X1 U181 ( .A(n102), .B(n53), .Y(P3[6]) );
  XNOR2X1 U182 ( .A(n102), .B(P13[9]), .Y(P2[0]) );
  XNOR2X1 U183 ( .A(n38), .B(P15[0]), .Y(P3[4]) );
  XNOR2X1 U184 ( .A(n25), .B(P14[8]), .Y(P3[12]) );
  XOR2X1 U185 ( .A(n96), .B(P2[1]), .Y(P15[12]) );
  XNOR2X1 U186 ( .A(n135), .B(P6[2]), .Y(P2[7]) );
  XNOR2X1 U187 ( .A(n39), .B(n64), .Y(n27) );
  XNOR2X1 U188 ( .A(n12), .B(n127), .Y(P13[9]) );
  XNOR2X1 U189 ( .A(n12), .B(n154), .Y(n63) );
  XNOR2X1 U190 ( .A(n150), .B(n120), .Y(n104) );
  XNOR2X1 U191 ( .A(n102), .B(n153), .Y(n155) );
  XNOR2X1 U192 ( .A(n94), .B(n104), .Y(P10[2]) );
  XNOR2X1 U193 ( .A(n12), .B(P1[1]), .Y(P13[7]) );
  XNOR2X1 U194 ( .A(n12), .B(n126), .Y(n71) );
  XNOR2X1 U195 ( .A(n37), .B(n38), .Y(n36) );
  XNOR2X1 U196 ( .A(n135), .B(n116), .Y(P3[8]) );
  XNOR2X1 U197 ( .A(n8), .B(n52), .Y(P4[8]) );
  XNOR2X1 U198 ( .A(n102), .B(n152), .Y(P10[9]) );
  XNOR2X1 U199 ( .A(n12), .B(n101), .Y(P14[3]) );
  XNOR2X1 U200 ( .A(n94), .B(n122), .Y(P14[7]) );
  XNOR2XL U201 ( .A(n25), .B(n119), .Y(P3[1]) );
  XNOR2X1 U202 ( .A(n39), .B(n40), .Y(n35) );
  BUFX3 U203 ( .A(P2[11]), .Y(P1[4]) );
  BUFX3 U204 ( .A(P9[0]), .Y(P8[6]) );
  BUFX3 U205 ( .A(P15[4]), .Y(P16[11]) );
  BUFX2 U206 ( .A(P3[0]), .Y(P2[6]) );
  BUFX3 U207 ( .A(P2[4]), .Y(P3[11]) );
  BUFX3 U208 ( .A(P6[12]), .Y(P5[5]) );
  BUFX3 U209 ( .A(P5[4]), .Y(P6[11]) );
  XNOR2XL U210 ( .A(n42), .B(n207), .Y(P1[10]) );
  XNOR2X1 U211 ( .A(n7), .B(n31), .Y(P11[7]) );
  XNOR2X1 U212 ( .A(P1[11]), .B(n80), .Y(P16[7]) );
  XNOR2X1 U213 ( .A(n9), .B(n62), .Y(n122) );
  XOR2X1 U214 ( .A(n62), .B(n63), .Y(P8[12]) );
  XNOR2X1 U215 ( .A(n39), .B(n90), .Y(P13[6]) );
  XNOR2X1 U216 ( .A(n10), .B(n71), .Y(P7[0]) );
  XNOR2X1 U217 ( .A(n10), .B(n153), .Y(P11[4]) );
  XNOR2X1 U218 ( .A(n6), .B(n152), .Y(P12[12]) );
  XNOR2X1 U219 ( .A(n6), .B(n31), .Y(P9[4]) );
  XNOR2X1 U220 ( .A(n102), .B(n88), .Y(P4[6]) );
  XOR2X1 U221 ( .A(n24), .B(n72), .Y(P7[12]) );
  XOR2X1 U222 ( .A(n50), .B(n88), .Y(P6[12]) );
  XNOR2XL U223 ( .A(n7), .B(b[8]), .Y(n134) );
  XNOR2XL U224 ( .A(n6), .B(b[9]), .Y(n89) );
  XNOR2X1 U225 ( .A(P6[2]), .B(n140), .Y(P8[5]) );
  XOR2X1 U226 ( .A(n12), .B(n207), .Y(n140) );
  XNOR2X1 U227 ( .A(n11), .B(n122), .Y(P12[1]) );
  XNOR2X1 U228 ( .A(n10), .B(n133), .Y(n116) );
  XNOR2X1 U229 ( .A(n30), .B(n139), .Y(P14[8]) );
  XNOR2XL U230 ( .A(n25), .B(n207), .Y(n85) );
  XNOR2X1 U231 ( .A(n7), .B(P7[1]), .Y(n53) );
  XOR2XL U232 ( .A(P1[11]), .B(P1[0]), .Y(n156) );
  XNOR2X1 U233 ( .A(n48), .B(n93), .Y(n120) );
  XOR2X1 U234 ( .A(n128), .B(P1[1]), .Y(n153) );
  XOR2X1 U235 ( .A(n59), .B(n147), .Y(n139) );
  XNOR2XL U236 ( .A(n70), .B(b[9]), .Y(n147) );
  XNOR2X1 U237 ( .A(n76), .B(n95), .Y(P16[1]) );
  XOR2X1 U238 ( .A(n109), .B(n72), .Y(P16[3]) );
  XNOR2X1 U239 ( .A(n9), .B(n114), .Y(n73) );
  XNOR2X1 U240 ( .A(n30), .B(n96), .Y(n154) );
  INVX1 U241 ( .A(P12[7]), .Y(n51) );
  XNOR2X1 U242 ( .A(n7), .B(n28), .Y(P6[2]) );
  XNOR2X1 U243 ( .A(b[4]), .B(n42), .Y(P12[8]) );
  XOR2X1 U244 ( .A(n58), .B(n62), .Y(n55) );
  XOR2X1 U245 ( .A(n157), .B(n40), .Y(n26) );
  XOR2X1 U246 ( .A(n5), .B(n207), .Y(n157) );
  XOR2X1 U247 ( .A(n68), .B(n69), .Y(n41) );
  XOR2X1 U248 ( .A(b[8]), .B(n85), .Y(n58) );
  INVX1 U249 ( .A(n86), .Y(n38) );
  XOR2X1 U250 ( .A(P14[2]), .B(n138), .Y(P15[10]) );
  XNOR2X1 U251 ( .A(n67), .B(n82), .Y(P5[8]) );
  XNOR2X1 U252 ( .A(n6), .B(n34), .Y(P9[2]) );
  XNOR2X1 U253 ( .A(n6), .B(n56), .Y(P12[10]) );
  XNOR2XL U254 ( .A(n135), .B(n136), .Y(P15[2]) );
  XNOR2X1 U255 ( .A(n9), .B(n53), .Y(P8[2]) );
  XNOR2X1 U256 ( .A(n7), .B(n101), .Y(P4[7]) );
  XNOR2X1 U257 ( .A(b[9]), .B(n99), .Y(P4[9]) );
  XOR2X1 U258 ( .A(n129), .B(n130), .Y(P15[9]) );
  XOR2X1 U259 ( .A(n90), .B(P13[10]), .Y(n130) );
  XOR2X1 U260 ( .A(n62), .B(n116), .Y(P11[2]) );
  BUFX3 U261 ( .A(P10[5]), .Y(P11[12]) );
  BUFX3 U262 ( .A(P11[4]), .Y(P12[11]) );
  BUFX3 U263 ( .A(P10[12]), .Y(P9[5]) );
  XOR2X1 U264 ( .A(n90), .B(n46), .Y(n79) );
  XNOR2X1 U265 ( .A(n118), .B(n135), .Y(n49) );
  XNOR2X1 U266 ( .A(b[9]), .B(n108), .Y(P16[6]) );
  XNOR2XL U267 ( .A(n135), .B(n117), .Y(P10[1]) );
  XNOR2X1 U268 ( .A(P11[7]), .B(n94), .Y(P5[2]) );
  XOR2X1 U269 ( .A(P1[2]), .B(n142), .Y(P14[1]) );
  BUFX3 U270 ( .A(P8[12]), .Y(P7[5]) );
  BUFX3 U271 ( .A(P4[12]), .Y(P3[5]) );
  BUFX3 U272 ( .A(P4[4]), .Y(P5[11]) );
  CLKBUFXL U273 ( .A(P12[4]), .Y(P13[11]) );
  BUFX3 U274 ( .A(P13[5]), .Y(P14[12]) );
  CLKBUFXL U275 ( .A(P7[4]), .Y(P8[11]) );
  XNOR2X1 U276 ( .A(n25), .B(n63), .Y(P11[1]) );
  XNOR2X1 U277 ( .A(n9), .B(n155), .Y(P11[10]) );
  XNOR2X1 U278 ( .A(b[11]), .B(n99), .Y(P10[3]) );
  XNOR2X1 U280 ( .A(n135), .B(n155), .Y(P10[8]) );
  BUFX3 U281 ( .A(P9[4]), .Y(P10[11]) );
  XNOR2X1 U282 ( .A(n7), .B(P2[11]), .Y(P8[9]) );
  BUFX3 U283 ( .A(P8[0]), .Y(P7[6]) );
  BUFX3 U284 ( .A(P4[6]), .Y(P5[0]) );
  XNOR2X1 U285 ( .A(b[11]), .B(n95), .Y(P5[1]) );
  XOR2X1 U286 ( .A(P11[7]), .B(n112), .Y(P4[1]) );
  BUFX3 U287 ( .A(P13[6]), .Y(P14[0]) );
  BUFX3 U288 ( .A(P7[0]), .Y(P6[6]) );
  BUFX3 U289 ( .A(P6[4]), .Y(P7[11]) );
  XNOR2X1 U290 ( .A(n67), .B(n41), .Y(P6[7]) );
  BUFX3 U291 ( .A(P8[5]), .Y(P9[12]) );
  BUFX3 U292 ( .A(P7[12]), .Y(P6[5]) );
  XNOR2X1 U293 ( .A(n83), .B(n82), .Y(P5[7]) );
  XOR2X1 U294 ( .A(n58), .B(n59), .Y(P7[7]) );
  XNOR2X1 U295 ( .A(n51), .B(n52), .Y(P8[3]) );
  XNOR2X1 U296 ( .A(P1[0]), .B(n78), .Y(P4[10]) );
  CLKBUFXL U297 ( .A(P13[0]), .Y(P12[6]) );
  XOR2X1 U298 ( .A(n96), .B(P7[3]), .Y(P5[10]) );
  XNOR2XL U299 ( .A(n207), .B(n111), .Y(P4[2]) );
  XNOR2X1 U300 ( .A(n39), .B(n139), .Y(P12[2]) );
  XOR2X1 U301 ( .A(n35), .B(n36), .Y(P9[1]) );
  XNOR2X1 U302 ( .A(n8), .B(n33), .Y(P9[3]) );
  BUFX3 U303 ( .A(P8[4]), .Y(P9[11]) );
  XOR2XL U304 ( .A(n62), .B(n117), .Y(P3[3]) );
  XNOR2X1 U305 ( .A(n25), .B(P7[2]), .Y(P3[7]) );
  XNOR2X1 U306 ( .A(n9), .B(n115), .Y(P3[9]) );
  XNOR2X1 U307 ( .A(n6), .B(n120), .Y(P3[10]) );
  BUFX3 U308 ( .A(P3[12]), .Y(P2[5]) );
  XNOR2X1 U309 ( .A(n10), .B(P13[10]), .Y(P1[7]) );
  BUFX3 U310 ( .A(P15[11]), .Y(P14[4]) );
  XNOR2X1 U311 ( .A(n115), .B(n37), .Y(n148) );
  XNOR2X1 U312 ( .A(n21), .B(n22), .Y(n20) );
  BUFX3 U313 ( .A(P12[12]), .Y(P11[5]) );
  XNOR2XL U314 ( .A(n135), .B(P1[0]), .Y(n112) );
  XOR2X1 U315 ( .A(b_0), .B(n154), .Y(n115) );
  XOR2X1 U316 ( .A(b_2), .B(n151), .Y(P12[0]) );
  XNOR2X1 U317 ( .A(n60), .B(n158), .Y(P8[0]) );
  XOR2XL U318 ( .A(b_3), .B(b[11]), .Y(n59) );
  XNOR2X2 U319 ( .A(b_3), .B(n39), .Y(n83) );
  XNOR2X1 U320 ( .A(b_2), .B(n57), .Y(n118) );
  XOR2X1 U321 ( .A(n73), .B(P1[10]), .Y(n146) );
  XNOR2X1 U322 ( .A(b_1), .B(n87), .Y(P16[4]) );
  XNOR2X1 U323 ( .A(n77), .B(n78), .Y(P6[3]) );
  XNOR2X1 U324 ( .A(n7), .B(n66), .Y(P6[8]) );
  XNOR2X1 U325 ( .A(n25), .B(b_0), .Y(n69) );
  XNOR2X1 U326 ( .A(n39), .B(b_0), .Y(n125) );
  XNOR2X1 U327 ( .A(n8), .B(P13[5]), .Y(P2[9]) );
  XNOR2X1 U328 ( .A(n3), .B(n79), .Y(P6[10]) );
  XNOR2X1 U329 ( .A(n3), .B(n26), .Y(P6[4]) );
  XNOR2X1 U330 ( .A(n3), .B(n59), .Y(n60) );
  XNOR2X1 U331 ( .A(b_3), .B(n3), .Y(P12[7]) );
  XNOR2X1 U332 ( .A(P1[11]), .B(n74), .Y(P13[2]) );
  XOR2X1 U333 ( .A(n67), .B(n143), .Y(P13[3]) );
  XNOR2X1 U334 ( .A(n39), .B(n67), .Y(n28) );
  XNOR2X1 U335 ( .A(n5), .B(n41), .Y(P9[10]) );
  XNOR2X1 U336 ( .A(n5), .B(n49), .Y(P3[2]) );
  XNOR2X1 U337 ( .A(n5), .B(n148), .Y(P11[9]) );
  XNOR2XL U338 ( .A(n7), .B(n5), .Y(n129) );
  XNOR2X1 U339 ( .A(n47), .B(n70), .Y(n92) );
  XOR2X1 U340 ( .A(n44), .B(P2[9]), .Y(P8[7]) );
  XNOR2X1 U341 ( .A(n11), .B(n60), .Y(P14[10]) );
  XNOR2X1 U342 ( .A(n11), .B(n24), .Y(P9[8]) );
  XNOR2X1 U343 ( .A(n11), .B(n71), .Y(P16[2]) );
  XNOR2X1 U344 ( .A(n11), .B(n125), .Y(n56) );
  XOR2X1 U345 ( .A(b[5]), .B(n207), .Y(n107) );
  XNOR2X1 U346 ( .A(n11), .B(n98), .Y(P7[1]) );
  XNOR2XL U347 ( .A(n23), .B(b[11]), .Y(n37) );
  XNOR2XL U348 ( .A(n11), .B(P1[0]), .Y(n141) );
  XOR2X1 U349 ( .A(b[5]), .B(b[8]), .Y(n90) );
  XNOR2X1 U350 ( .A(b[5]), .B(n74), .Y(n67) );
  XNOR2X1 U351 ( .A(n54), .B(b_2), .Y(n93) );
  XNOR2X1 U352 ( .A(n54), .B(n77), .Y(P13[5]) );
  XNOR2X1 U353 ( .A(n102), .B(n19), .Y(P13[10]) );
  XOR2X1 U354 ( .A(n19), .B(n20), .Y(P9[9]) );
  XOR2X1 U355 ( .A(P2[2]), .B(n93), .Y(P5[3]) );
  XNOR2X1 U356 ( .A(n1), .B(n106), .Y(P4[5]) );
  XOR2X1 U357 ( .A(P1[5]), .B(n141), .Y(n101) );
  XNOR2XL U358 ( .A(n12), .B(n149), .Y(P11[0]) );
  XNOR2X1 U359 ( .A(n13), .B(n121), .Y(P14[9]) );
  XNOR2X1 U360 ( .A(n13), .B(n56), .Y(P7[9]) );
  XNOR2X1 U361 ( .A(b[10]), .B(n148), .Y(P10[7]) );
  XNOR2X1 U362 ( .A(n13), .B(P6[1]), .Y(P3[0]) );
  XNOR2X1 U363 ( .A(n13), .B(n151), .Y(P10[5]) );
  XNOR2X1 U364 ( .A(n13), .B(n46), .Y(P9[0]) );
  XNOR2X1 U365 ( .A(n13), .B(n96), .Y(P7[2]) );
  XNOR2X1 U366 ( .A(n13), .B(P13[7]), .Y(P2[11]) );
  XNOR2X2 U367 ( .A(b_3), .B(n45), .Y(n86) );
endmodule


module multiplier_column6_p16 ( b, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, 
        P11, P12, P13, P14, P15, P16 );
  input [12:0] b;
  output [12:0] P1;
  output [12:0] P2;
  output [12:0] P3;
  output [12:0] P4;
  output [12:0] P5;
  output [12:0] P6;
  output [12:0] P7;
  output [12:0] P8;
  output [12:0] P9;
  output [12:0] P10;
  output [12:0] P11;
  output [12:0] P12;
  output [12:0] P13;
  output [12:0] P14;
  output [12:0] P15;
  output [12:0] P16;
  wire   b_3, b_2, b_1, b_0, n253, n18, n19, n20, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n38, n39, n40, n41, n42,
         n44, n45, n46, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n127,
         n128, n129, n130, n131, n132, n133, n1, n2, n3, n4, n5, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n21, n37, n43, n47, n48, n65, n78,
         n81, n109, n126, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n212, n213, n215, n216,
         n217, n218;
  assign b_3 = b[3];
  assign b_2 = b[2];
  assign b_1 = b[1];
  assign b_0 = b[0];

  CLKINVX2 U1 ( .A(b[8]), .Y(n47) );
  XNOR2X4 U2 ( .A(n97), .B(b[7]), .Y(n25) );
  CLKINVX3 U3 ( .A(n213), .Y(n58) );
  XNOR2X2 U4 ( .A(n218), .B(n25), .Y(P15[4]) );
  CLKBUFXL U5 ( .A(n253), .Y(P16[3]) );
  XNOR2X1 U6 ( .A(n17), .B(n88), .Y(n101) );
  XNOR2X2 U7 ( .A(n213), .B(n49), .Y(n110) );
  NAND2X1 U8 ( .A(n134), .B(n135), .Y(P14[6]) );
  NAND2BXL U9 ( .AN(b[6]), .B(n52), .Y(n15) );
  OAI21XL U10 ( .A0(n94), .A1(n84), .B0(n136), .Y(P4[2]) );
  OAI2BB1X2 U11 ( .A0N(n215), .A1N(n37), .B0(n43), .Y(P3[0]) );
  INVX1 U12 ( .A(P15[4]), .Y(n37) );
  XNOR2XL U13 ( .A(n218), .B(b[9]), .Y(n131) );
  XNOR2XL U14 ( .A(n44), .B(n82), .Y(P13[2]) );
  XNOR2X4 U15 ( .A(b_2), .B(n22), .Y(n107) );
  INVX8 U16 ( .A(n215), .Y(n22) );
  CLKINVX3 U17 ( .A(n212), .Y(n32) );
  XNOR2X1 U18 ( .A(P3[0]), .B(n213), .Y(n24) );
  NAND2X2 U19 ( .A(n8), .B(n9), .Y(n11) );
  INVX1 U20 ( .A(n74), .Y(n8) );
  NAND2X2 U21 ( .A(n14), .B(n15), .Y(P4[6]) );
  INVX1 U22 ( .A(n52), .Y(n13) );
  XOR2X2 U23 ( .A(n216), .B(P15[8]), .Y(P2[11]) );
  XNOR2X2 U24 ( .A(n45), .B(n107), .Y(n89) );
  XOR2X1 U25 ( .A(n109), .B(n212), .Y(n146) );
  XNOR2XL U26 ( .A(n3), .B(n104), .Y(P16[9]) );
  XOR2X1 U27 ( .A(n213), .B(n104), .Y(n82) );
  XNOR2XL U28 ( .A(n218), .B(n101), .Y(n27) );
  INVX1 U29 ( .A(n17), .Y(n21) );
  XOR2X1 U30 ( .A(P1[9]), .B(P2[0]), .Y(n87) );
  XNOR2X1 U31 ( .A(n124), .B(n1), .Y(n20) );
  CLKINVX3 U32 ( .A(b[4]), .Y(n97) );
  XNOR2X1 U33 ( .A(P1[10]), .B(P14[4]), .Y(n124) );
  BUFX3 U34 ( .A(b[8]), .Y(n215) );
  INVX1 U35 ( .A(b_1), .Y(n109) );
  XNOR2X1 U36 ( .A(n34), .B(n64), .Y(n104) );
  BUFX3 U37 ( .A(P3[0]), .Y(P2[7]) );
  CLKINVX3 U38 ( .A(b[11]), .Y(n29) );
  BUFX3 U39 ( .A(b[5]), .Y(P1[11]) );
  XNOR2X1 U40 ( .A(n63), .B(n83), .Y(n33) );
  NAND2X1 U41 ( .A(n134), .B(n135), .Y(P15[12]) );
  INVX1 U42 ( .A(n110), .Y(n126) );
  NAND2X1 U43 ( .A(b[6]), .B(n13), .Y(n14) );
  CLKINVX3 U44 ( .A(b[9]), .Y(n44) );
  INVX2 U45 ( .A(b[12]), .Y(n34) );
  XOR2X2 U46 ( .A(n88), .B(n89), .Y(n52) );
  XNOR2X1 U47 ( .A(n119), .B(n29), .Y(P8[9]) );
  XNOR2X1 U48 ( .A(n58), .B(n94), .Y(P2[0]) );
  XNOR2X2 U49 ( .A(P2[11]), .B(n212), .Y(n18) );
  CLKBUFX8 U50 ( .A(b_0), .Y(n212) );
  XNOR2XL U51 ( .A(n95), .B(P1[10]), .Y(n84) );
  XNOR2XL U52 ( .A(n22), .B(P1[10]), .Y(n142) );
  XOR2X1 U53 ( .A(P1[10]), .B(P8[1]), .Y(P4[10]) );
  BUFX3 U54 ( .A(b[4]), .Y(P1[10]) );
  INVX1 U55 ( .A(b[7]), .Y(n1) );
  XNOR2XL U56 ( .A(n12), .B(P15[1]), .Y(n80) );
  XNOR2X1 U57 ( .A(n63), .B(n100), .Y(P8[1]) );
  INVX1 U58 ( .A(b[6]), .Y(n63) );
  INVX1 U59 ( .A(b_3), .Y(n3) );
  INVX1 U60 ( .A(b_3), .Y(n2) );
  INVX1 U61 ( .A(b_2), .Y(n4) );
  XNOR2X1 U62 ( .A(n4), .B(n127), .Y(P11[8]) );
  XNOR2XL U63 ( .A(n4), .B(b[10]), .Y(n61) );
  XNOR2X1 U64 ( .A(n117), .B(n4), .Y(P13[7]) );
  INVX1 U65 ( .A(b_2), .Y(n49) );
  INVX1 U66 ( .A(P1[11]), .Y(n5) );
  XNOR2XL U67 ( .A(n31), .B(n218), .Y(n75) );
  XNOR2X1 U68 ( .A(n124), .B(n218), .Y(n115) );
  XNOR2XL U69 ( .A(b_2), .B(n218), .Y(n54) );
  XNOR2X2 U70 ( .A(n218), .B(n212), .Y(n111) );
  XOR2XL U71 ( .A(n216), .B(n213), .Y(n144) );
  XNOR2XL U72 ( .A(n216), .B(n1), .Y(n91) );
  XNOR2XL U73 ( .A(n216), .B(n49), .Y(n112) );
  XOR2XL U74 ( .A(n216), .B(b[11]), .Y(n69) );
  BUFX3 U75 ( .A(b[12]), .Y(n216) );
  BUFX3 U76 ( .A(b[7]), .Y(P1[0]) );
  XNOR2X1 U77 ( .A(P1[0]), .B(n39), .Y(P7[9]) );
  XOR2X1 U78 ( .A(n32), .B(P1[0]), .Y(n141) );
  XNOR2XL U79 ( .A(n22), .B(P1[0]), .Y(P1[1]) );
  XNOR2X1 U80 ( .A(b_2), .B(P1[0]), .Y(n74) );
  INVX1 U81 ( .A(b[7]), .Y(n72) );
  XNOR2X4 U82 ( .A(n29), .B(P1[2]), .Y(P15[8]) );
  BUFX1 U83 ( .A(n97), .Y(n217) );
  NAND2X1 U84 ( .A(n74), .B(P15[2]), .Y(n10) );
  NAND2X4 U85 ( .A(n10), .B(n11), .Y(n133) );
  INVX2 U86 ( .A(P15[2]), .Y(n9) );
  XNOR2X2 U87 ( .A(n3), .B(n111), .Y(P15[2]) );
  INVX1 U88 ( .A(b[6]), .Y(n12) );
  XNOR2X4 U89 ( .A(P4[6]), .B(n79), .Y(n59) );
  DLY1X1 U90 ( .A(P4[6]), .Y(P5[12]) );
  XNOR2XL U91 ( .A(n44), .B(n100), .Y(P15[9]) );
  INVXL U92 ( .A(n64), .Y(n17) );
  XOR2X1 U93 ( .A(b[10]), .B(b[11]), .Y(n94) );
  XNOR2X1 U94 ( .A(n82), .B(b[5]), .Y(n16) );
  XNOR2XL U95 ( .A(n82), .B(b[5]), .Y(n41) );
  NAND2XL U96 ( .A(n47), .B(P15[4]), .Y(n43) );
  NAND2X1 U97 ( .A(n48), .B(n65), .Y(n81) );
  NAND2X1 U98 ( .A(n78), .B(n81), .Y(n253) );
  INVX1 U99 ( .A(n71), .Y(n65) );
  XNOR2X1 U100 ( .A(n49), .B(b_3), .Y(P15[0]) );
  XNOR2X1 U101 ( .A(b[10]), .B(n1), .Y(n71) );
  NAND2XL U102 ( .A(n18), .B(n71), .Y(n78) );
  INVX1 U103 ( .A(n18), .Y(n48) );
  XOR2X1 U104 ( .A(P1[0]), .B(n120), .Y(n119) );
  XNOR2X2 U105 ( .A(b[10]), .B(n34), .Y(n100) );
  BUFX3 U106 ( .A(P8[12]), .Y(P7[6]) );
  XNOR2X1 U107 ( .A(n217), .B(P2[1]), .Y(P16[7]) );
  XNOR2X1 U108 ( .A(n217), .B(n87), .Y(P2[3]) );
  BUFX3 U109 ( .A(P5[4]), .Y(P6[10]) );
  XNOR2X1 U110 ( .A(n217), .B(n111), .Y(P14[9]) );
  XNOR2X1 U111 ( .A(n22), .B(n216), .Y(n138) );
  XNOR2X1 U112 ( .A(n5), .B(n120), .Y(P13[4]) );
  XOR2XL U113 ( .A(n58), .B(P1[0]), .Y(n145) );
  XNOR2XL U114 ( .A(n4), .B(n129), .Y(P12[1]) );
  XOR2X1 U115 ( .A(P8[5]), .B(n70), .Y(P6[1]) );
  XNOR2X1 U116 ( .A(b_3), .B(n1), .Y(n85) );
  XOR2XL U117 ( .A(n29), .B(b[5]), .Y(n149) );
  NAND2XL U118 ( .A(n34), .B(n110), .Y(n134) );
  NAND2X1 U119 ( .A(b[12]), .B(n126), .Y(n135) );
  NAND2XL U120 ( .A(n94), .B(n84), .Y(n136) );
  XOR2XL U121 ( .A(n4), .B(n212), .Y(n148) );
  XOR2XL U122 ( .A(n4), .B(b[9]), .Y(n143) );
  CLKBUFXL U123 ( .A(P13[10]), .Y(P12[4]) );
  XNOR2XL U124 ( .A(n1), .B(n98), .Y(P3[7]) );
  BUFX2 U125 ( .A(P11[11]), .Y(P10[5]) );
  CLKBUFXL U126 ( .A(P15[4]), .Y(P16[10]) );
  CLKBUFXL U127 ( .A(P12[5]), .Y(P13[11]) );
  CLKBUFXL U128 ( .A(P2[0]), .Y(P1[7]) );
  XNOR2XL U129 ( .A(n12), .B(n86), .Y(P16[12]) );
  XOR2XL U130 ( .A(n137), .B(n21), .Y(n92) );
  XNOR2XL U131 ( .A(n212), .B(P15[8]), .Y(n137) );
  XNOR2XL U132 ( .A(n32), .B(n88), .Y(n106) );
  XOR2X1 U133 ( .A(n94), .B(n138), .Y(P16[2]) );
  XOR2X1 U134 ( .A(b[11]), .B(n33), .Y(n127) );
  XOR2X1 U135 ( .A(n139), .B(n70), .Y(n99) );
  XOR2XL U136 ( .A(n216), .B(n212), .Y(n139) );
  XNOR2XL U137 ( .A(n218), .B(P1[10]), .Y(n53) );
  XNOR2X1 U138 ( .A(n140), .B(n30), .Y(n90) );
  XNOR2XL U139 ( .A(n216), .B(b[9]), .Y(n140) );
  XNOR2XL U140 ( .A(n2), .B(P1[10]), .Y(P14[8]) );
  XNOR2XL U141 ( .A(n12), .B(n99), .Y(P3[6]) );
  XNOR2XL U142 ( .A(n5), .B(n95), .Y(P11[11]) );
  XNOR2X1 U143 ( .A(P8[3]), .B(n141), .Y(P6[12]) );
  XNOR2X1 U144 ( .A(n36), .B(n142), .Y(P9[12]) );
  XNOR2X1 U145 ( .A(n26), .B(n143), .Y(P11[12]) );
  XNOR2X1 U146 ( .A(n59), .B(n144), .Y(P5[4]) );
  CLKBUFXL U147 ( .A(P2[11]), .Y(P1[5]) );
  XNOR2X4 U148 ( .A(n47), .B(b[9]), .Y(P1[2]) );
  XNOR2X1 U149 ( .A(b[11]), .B(n44), .Y(n88) );
  XNOR2XL U150 ( .A(n58), .B(P1[10]), .Y(n57) );
  XNOR2X1 U151 ( .A(n83), .B(n145), .Y(n30) );
  XOR2X1 U152 ( .A(n63), .B(n146), .Y(n120) );
  XNOR2XL U153 ( .A(n12), .B(n46), .Y(P15[3]) );
  XNOR2XL U154 ( .A(n212), .B(n31), .Y(P9[1]) );
  XOR2XL U155 ( .A(n56), .B(n55), .Y(P6[8]) );
  XNOR2X1 U156 ( .A(n29), .B(n30), .Y(P9[2]) );
  CLKBUFXL U157 ( .A(P4[10]), .Y(P3[4]) );
  CLKBUFXL U158 ( .A(P5[0]), .Y(P4[7]) );
  XNOR2XL U159 ( .A(n3), .B(n23), .Y(P10[9]) );
  CLKBUFXL U160 ( .A(P15[0]), .Y(P14[7]) );
  CLKBUFXL U161 ( .A(P14[4]), .Y(P15[10]) );
  XOR2X1 U162 ( .A(n60), .B(n62), .Y(P6[5]) );
  XNOR2XL U163 ( .A(n2), .B(n212), .Y(n62) );
  XNOR2X1 U164 ( .A(b_2), .B(n217), .Y(P15[1]) );
  XNOR2X1 U165 ( .A(b[6]), .B(n97), .Y(n64) );
  XOR2X1 U166 ( .A(n147), .B(n131), .Y(n23) );
  XOR2X1 U167 ( .A(b[6]), .B(n112), .Y(n147) );
  XNOR2XL U168 ( .A(b[6]), .B(P1[0]), .Y(n132) );
  XOR2X1 U169 ( .A(n60), .B(n61), .Y(P7[12]) );
  BUFX8 U170 ( .A(n76), .Y(n218) );
  CLKBUFXL U171 ( .A(b[6]), .Y(P1[12]) );
  XNOR2X1 U172 ( .A(P8[9]), .B(n77), .Y(P13[10]) );
  BUFX3 U173 ( .A(P11[5]), .Y(P12[11]) );
  BUFX3 U174 ( .A(P12[12]), .Y(P11[6]) );
  BUFX3 U175 ( .A(P12[0]), .Y(P11[7]) );
  BUFX3 U176 ( .A(P13[12]), .Y(P12[6]) );
  BUFX3 U177 ( .A(P2[12]), .Y(P1[6]) );
  BUFX3 U178 ( .A(P3[12]), .Y(P2[6]) );
  BUFX3 U179 ( .A(P6[0]), .Y(P5[7]) );
  BUFX3 U180 ( .A(P5[10]), .Y(P4[4]) );
  BUFX3 U181 ( .A(P10[4]), .Y(P11[10]) );
  BUFX3 U182 ( .A(P8[4]), .Y(P9[10]) );
  BUFX3 U183 ( .A(P9[4]), .Y(P10[10]) );
  XOR2X1 U184 ( .A(n86), .B(n87), .Y(P5[0]) );
  XOR2X1 U185 ( .A(P15[12]), .B(n53), .Y(P7[1]) );
  XNOR2X1 U186 ( .A(n29), .B(n130), .Y(n114) );
  XNOR2X1 U187 ( .A(n44), .B(n110), .Y(n98) );
  XNOR2X1 U188 ( .A(n58), .B(n69), .Y(n108) );
  XNOR2X1 U189 ( .A(n68), .B(n123), .Y(n93) );
  XNOR2X1 U190 ( .A(n217), .B(n131), .Y(n35) );
  XNOR2X1 U191 ( .A(n1), .B(n99), .Y(n51) );
  XOR2X1 U192 ( .A(n110), .B(P14[8]), .Y(n46) );
  XNOR2X1 U193 ( .A(n32), .B(n108), .Y(P15[11]) );
  XNOR2X1 U194 ( .A(n32), .B(n117), .Y(P12[12]) );
  XNOR2X1 U195 ( .A(n32), .B(P15[9]), .Y(P2[12]) );
  XNOR2X1 U196 ( .A(n29), .B(P7[2]), .Y(P2[5]) );
  XNOR2X1 U197 ( .A(n29), .B(P15[7]), .Y(P2[10]) );
  XNOR2X1 U198 ( .A(n44), .B(n118), .Y(P13[12]) );
  XNOR2X1 U199 ( .A(n44), .B(n42), .Y(P8[12]) );
  XNOR2X1 U200 ( .A(n58), .B(n116), .Y(P12[0]) );
  XNOR2X1 U201 ( .A(n58), .B(n118), .Y(P14[12]) );
  XNOR2X1 U202 ( .A(P11[2]), .B(n77), .Y(P6[0]) );
  XNOR2X1 U203 ( .A(n91), .B(n92), .Y(P5[10]) );
  XNOR2X1 U204 ( .A(n217), .B(n51), .Y(P10[4]) );
  XNOR2X1 U205 ( .A(n72), .B(P16[9]), .Y(P3[12]) );
  XNOR2X1 U206 ( .A(n34), .B(n118), .Y(P11[5]) );
  XNOR2X1 U207 ( .A(n34), .B(n35), .Y(P9[0]) );
  XOR2X1 U208 ( .A(P2[1]), .B(n38), .Y(P8[4]) );
  XOR2X1 U209 ( .A(n25), .B(n26), .Y(P9[4]) );
  XNOR2X1 U210 ( .A(n36), .B(n131), .Y(P4[9]) );
  XNOR2X1 U211 ( .A(n1), .B(n40), .Y(P8[2]) );
  XOR2X1 U212 ( .A(n32), .B(P2[0]), .Y(n68) );
  XNOR2X1 U213 ( .A(n29), .B(P1[3]), .Y(P16[1]) );
  XNOR2XL U214 ( .A(n34), .B(n89), .Y(P16[5]) );
  XNOR2X1 U215 ( .A(n24), .B(n38), .Y(n60) );
  BUFX3 U216 ( .A(P11[4]), .Y(P12[10]) );
  BUFX3 U217 ( .A(P14[11]), .Y(P13[5]) );
  XOR2X1 U218 ( .A(n91), .B(n114), .Y(P11[9]) );
  XNOR2X1 U219 ( .A(n217), .B(P16[12]), .Y(P3[1]) );
  XNOR2X1 U220 ( .A(n217), .B(P16[6]), .Y(P3[9]) );
  XNOR2X1 U221 ( .A(n1), .B(n102), .Y(P3[2]) );
  XNOR2X1 U222 ( .A(n1), .B(n27), .Y(P3[3]) );
  XNOR2X1 U223 ( .A(n112), .B(n96), .Y(P14[3]) );
  XNOR2X1 U224 ( .A(n27), .B(n28), .Y(P9[3]) );
  XOR2X1 U225 ( .A(n69), .B(P13[7]), .Y(P6[2]) );
  XOR2X1 U226 ( .A(P7[1]), .B(n122), .Y(P10[8]) );
  XOR2X1 U227 ( .A(P15[2]), .B(n122), .Y(P13[1]) );
  BUFX3 U228 ( .A(P6[4]), .Y(P7[10]) );
  BUFX3 U229 ( .A(P15[7]), .Y(P16[0]) );
  BUFX3 U230 ( .A(P13[7]), .Y(P14[0]) );
  BUFX3 U231 ( .A(P8[5]), .Y(P9[11]) );
  BUFX3 U232 ( .A(P10[0]), .Y(P9[7]) );
  BUFX3 U233 ( .A(P9[5]), .Y(P10[11]) );
  BUFX3 U234 ( .A(P7[0]), .Y(P6[7]) );
  BUFX3 U235 ( .A(P13[0]), .Y(P12[7]) );
  BUFX3 U236 ( .A(P7[5]), .Y(P8[11]) );
  BUFX3 U237 ( .A(P2[4]), .Y(P3[10]) );
  BUFX3 U238 ( .A(P13[4]), .Y(P14[10]) );
  BUFX3 U239 ( .A(P6[5]), .Y(P7[11]) );
  BUFX3 U240 ( .A(P11[12]), .Y(P10[6]) );
  BUFX3 U241 ( .A(P11[0]), .Y(P10[7]) );
  BUFX3 U242 ( .A(P6[12]), .Y(P5[6]) );
  XOR2X1 U243 ( .A(n86), .B(n108), .Y(P16[4]) );
  INVX1 U244 ( .A(n123), .Y(n77) );
  BUFX3 U245 ( .A(P15[5]), .Y(P16[11]) );
  XOR2X1 U246 ( .A(n21), .B(n66), .Y(P6[4]) );
  XOR2X1 U247 ( .A(P1[10]), .B(n113), .Y(n117) );
  XNOR2X1 U248 ( .A(b[9]), .B(n72), .Y(n86) );
  XNOR2X1 U249 ( .A(n28), .B(n85), .Y(n118) );
  XNOR2X1 U250 ( .A(n32), .B(n94), .Y(P14[4]) );
  XNOR2X1 U251 ( .A(n218), .B(n67), .Y(P15[5]) );
  XNOR2X1 U252 ( .A(n29), .B(P15[0]), .Y(P2[2]) );
  XNOR2X1 U253 ( .A(n103), .B(P1[1]), .Y(P15[7]) );
  XOR2X1 U254 ( .A(n71), .B(P2[2]), .Y(P8[5]) );
  XNOR2X1 U255 ( .A(n105), .B(n106), .Y(P16[6]) );
  XNOR2X1 U256 ( .A(n103), .B(P15[12]), .Y(P2[1]) );
  XNOR2X1 U257 ( .A(n103), .B(n86), .Y(P1[3]) );
  XNOR2X1 U258 ( .A(n50), .B(n71), .Y(n96) );
  XNOR2XL U259 ( .A(n12), .B(b[9]), .Y(n38) );
  XNOR2XL U260 ( .A(n58), .B(n215), .Y(n70) );
  XNOR2X1 U261 ( .A(n66), .B(b[9]), .Y(n121) );
  XNOR2X1 U262 ( .A(n32), .B(n56), .Y(n130) );
  XNOR2X1 U263 ( .A(n103), .B(n35), .Y(n116) );
  XOR2X1 U264 ( .A(n127), .B(n128), .Y(n73) );
  XNOR2XL U265 ( .A(n216), .B(n218), .Y(n123) );
  XNOR2X1 U266 ( .A(n4), .B(n51), .Y(P7[4]) );
  XNOR2X1 U267 ( .A(n4), .B(n119), .Y(P14[11]) );
  XNOR2X1 U268 ( .A(n3), .B(P2[9]), .Y(P10[0]) );
  XNOR2X1 U269 ( .A(n103), .B(P7[1]), .Y(P2[4]) );
  XNOR2X1 U270 ( .A(n103), .B(n117), .Y(P13[0]) );
  XNOR2X1 U271 ( .A(b[11]), .B(n24), .Y(P9[5]) );
  XNOR2X1 U272 ( .A(n215), .B(n125), .Y(P12[5]) );
  XNOR2X1 U273 ( .A(b[11]), .B(n125), .Y(P11[4]) );
  XNOR2X1 U274 ( .A(P1[0]), .B(n59), .Y(P7[0]) );
  XNOR2X1 U275 ( .A(n5), .B(P8[2]), .Y(P3[5]) );
  XOR2X1 U276 ( .A(P5[0]), .B(n80), .Y(P5[5]) );
  XOR2X1 U277 ( .A(n20), .B(n105), .Y(P11[0]) );
  XNOR2X1 U278 ( .A(n103), .B(n130), .Y(n26) );
  XNOR2X1 U279 ( .A(n45), .B(n46), .Y(n42) );
  XOR2X1 U280 ( .A(n213), .B(n101), .Y(n129) );
  XNOR2XL U281 ( .A(n12), .B(n215), .Y(n67) );
  XNOR2XL U282 ( .A(P4[10]), .B(b[9]), .Y(n31) );
  XNOR2X1 U283 ( .A(P1[3]), .B(n12), .Y(P2[9]) );
  XOR2X1 U284 ( .A(P15[1]), .B(P16[2]), .Y(P4[8]) );
  XOR2X1 U285 ( .A(n215), .B(n98), .Y(n95) );
  XOR2X1 U286 ( .A(n54), .B(n56), .Y(P7[2]) );
  XNOR2X1 U287 ( .A(n5), .B(P2[2]), .Y(P16[8]) );
  XOR2X1 U288 ( .A(n79), .B(P4[8]), .Y(P8[3]) );
  XNOR2X1 U289 ( .A(b[11]), .B(n32), .Y(n40) );
  XOR2XL U290 ( .A(n54), .B(n55), .Y(P6[9]) );
  XNOR2X1 U291 ( .A(n216), .B(n3), .Y(P1[9]) );
  XOR2X1 U292 ( .A(n3), .B(n69), .Y(n36) );
  XOR2X1 U293 ( .A(n129), .B(n128), .Y(P11[2]) );
  XOR2X1 U294 ( .A(n253), .B(n57), .Y(n55) );
  XOR2X1 U295 ( .A(n110), .B(P4[9]), .Y(P11[3]) );
  INVXL U296 ( .A(n107), .Y(n28) );
  XOR2X1 U297 ( .A(n16), .B(P15[0]), .Y(n39) );
  XOR2X1 U298 ( .A(n83), .B(P13[7]), .Y(P5[2]) );
  XNOR2X1 U299 ( .A(n50), .B(n148), .Y(P7[5]) );
  BUFX3 U300 ( .A(P9[0]), .Y(P8[7]) );
  XNOR2X1 U301 ( .A(n2), .B(n116), .Y(P13[8]) );
  XNOR2X1 U302 ( .A(n44), .B(n114), .Y(P14[2]) );
  XNOR2X1 U303 ( .A(n4), .B(n102), .Y(P14[1]) );
  XNOR2X1 U304 ( .A(n12), .B(n93), .Y(P12[9]) );
  XNOR2X1 U305 ( .A(b[11]), .B(n121), .Y(P10[3]) );
  XNOR2X1 U306 ( .A(n215), .B(n20), .Y(P9[8]) );
  XNOR2X1 U307 ( .A(P1[10]), .B(n121), .Y(P13[3]) );
  XNOR2X1 U308 ( .A(n212), .B(n96), .Y(P4[1]) );
  XNOR2X1 U309 ( .A(n84), .B(n85), .Y(P5[1]) );
  BUFX3 U310 ( .A(P5[11]), .Y(P4[5]) );
  BUFX3 U311 ( .A(P16[12]), .Y(P15[6]) );
  XNOR2X1 U312 ( .A(n44), .B(n73), .Y(P12[3]) );
  BUFX3 U313 ( .A(P7[4]), .Y(P8[10]) );
  XNOR2X1 U314 ( .A(n67), .B(n68), .Y(P6[3]) );
  BUFX3 U315 ( .A(P5[5]), .Y(P6[11]) );
  BUFX3 U316 ( .A(P3[7]), .Y(P4[0]) );
  BUFX3 U317 ( .A(P3[5]), .Y(P4[11]) );
  BUFX3 U318 ( .A(P3[6]), .Y(P4[12]) );
  BUFX3 U319 ( .A(P2[5]), .Y(P3[11]) );
  BUFX3 U320 ( .A(P9[12]), .Y(P8[6]) );
  BUFX3 U321 ( .A(P10[12]), .Y(P9[6]) );
  XOR2X1 U322 ( .A(n74), .B(n75), .Y(P5[8]) );
  XNOR2X1 U323 ( .A(n1), .B(n73), .Y(P5[9]) );
  XNOR2X1 U324 ( .A(b[9]), .B(n115), .Y(P12[8]) );
  XNOR2X1 U325 ( .A(n217), .B(n90), .Y(P10[2]) );
  XNOR2X1 U326 ( .A(n32), .B(n33), .Y(P8[8]) );
  XOR2X1 U327 ( .A(n52), .B(n53), .Y(P7[3]) );
  XNOR2XL U328 ( .A(n2), .B(n89), .Y(P3[8]) );
  XNOR2X1 U329 ( .A(n44), .B(P15[5]), .Y(P2[8]) );
  BUFX3 U330 ( .A(P2[10]), .Y(P1[4]) );
  XNOR2X1 U331 ( .A(n4), .B(n69), .Y(P1[8]) );
  BUFX3 U332 ( .A(P15[11]), .Y(P14[5]) );
  BUFX3 U333 ( .A(P14[12]), .Y(P13[6]) );
  XOR2X1 U334 ( .A(n85), .B(n93), .Y(P4[3]) );
  BUFX3 U335 ( .A(P7[12]), .Y(P6[6]) );
  BUFX3 U336 ( .A(P8[0]), .Y(P7[7]) );
  XNOR2XL U337 ( .A(n29), .B(n215), .Y(n122) );
  XNOR2X1 U338 ( .A(n63), .B(b_3), .Y(n56) );
  INVXL U339 ( .A(b[10]), .Y(n103) );
  XOR2X1 U340 ( .A(n132), .B(P15[12]), .Y(n125) );
  XNOR2X1 U341 ( .A(n42), .B(n149), .Y(P8[0]) );
  XNOR2X1 U342 ( .A(b[10]), .B(b_0), .Y(n45) );
  INVX2 U343 ( .A(b[5]), .Y(n76) );
  XNOR2X1 U344 ( .A(b_3), .B(n92), .Y(P10[1]) );
  XNOR2X1 U345 ( .A(b[6]), .B(n115), .Y(P13[9]) );
  BUFX3 U346 ( .A(b_1), .Y(n213) );
  XOR2X1 U347 ( .A(n18), .B(n19), .Y(P9[9]) );
  XNOR2X1 U348 ( .A(n213), .B(b_3), .Y(n105) );
  XOR2X1 U349 ( .A(n213), .B(n113), .Y(n50) );
  XNOR2X1 U350 ( .A(P1[0]), .B(n41), .Y(P5[3]) );
  XNOR2X1 U351 ( .A(n40), .B(n39), .Y(P7[8]) );
  XNOR2X1 U352 ( .A(P1[2]), .B(n2), .Y(n113) );
  XNOR2XL U353 ( .A(n213), .B(b[5]), .Y(n19) );
  XOR2X1 U354 ( .A(n100), .B(n133), .Y(P12[2]) );
  XOR2X2 U355 ( .A(n215), .B(n133), .Y(n66) );
  XNOR2X1 U356 ( .A(b[5]), .B(n2), .Y(n79) );
  XOR2X1 U357 ( .A(b[10]), .B(b[5]), .Y(n83) );
  XNOR2X1 U358 ( .A(n22), .B(P12[2]), .Y(P11[1]) );
  XNOR2X1 U359 ( .A(n22), .B(n90), .Y(P5[11]) );
  XNOR2X1 U360 ( .A(n22), .B(n23), .Y(P10[12]) );
  XNOR2X1 U361 ( .A(n22), .B(n83), .Y(n102) );
  XNOR2X1 U362 ( .A(n22), .B(b_3), .Y(n128) );
endmodule


module multiplier_column5_p16 ( b, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, 
        P11, P12, P13, P14, P15, P16 );
  input [12:0] b;
  output [12:0] P1;
  output [12:0] P2;
  output [12:0] P3;
  output [12:0] P4;
  output [12:0] P5;
  output [12:0] P6;
  output [12:0] P7;
  output [12:0] P8;
  output [12:0] P9;
  output [12:0] P10;
  output [12:0] P11;
  output [12:0] P12;
  output [12:0] P13;
  output [12:0] P14;
  output [12:0] P15;
  output [12:0] P16;
  wire   b_3, b_2, b_1, b_0, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n39,
         n40, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n67, n68, n69,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n108, n110, n112, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n124, n125, n126, n127,
         n128, n129, n131, n132, n133, n1, n2, n3, n4, n5, n6, n8, n9, n10,
         n11, n12, n13, n25, n38, n41, n66, n70, n82, n106, n107, n109, n111,
         n113, n211;
  assign b_3 = b[3];
  assign b_2 = b[2];
  assign b_1 = b[1];
  assign b_0 = b[0];

  INVX4 U1 ( .A(b_2), .Y(n16) );
  XOR2X2 U2 ( .A(n124), .B(n131), .Y(n64) );
  XNOR2XL U3 ( .A(n83), .B(n33), .Y(P10[1]) );
  XOR2X2 U4 ( .A(P1[10]), .B(b[12]), .Y(n53) );
  BUFX12 U5 ( .A(b[5]), .Y(P1[10]) );
  INVX1 U6 ( .A(b[9]), .Y(n9) );
  XNOR2X2 U7 ( .A(n16), .B(b[9]), .Y(n34) );
  XOR2X1 U8 ( .A(P3[3]), .B(n40), .Y(n37) );
  XNOR2XL U9 ( .A(n28), .B(P1[11]), .Y(n27) );
  XOR2X1 U10 ( .A(n32), .B(n33), .Y(P8[5]) );
  XNOR2X1 U11 ( .A(n52), .B(b[7]), .Y(n36) );
  INVX2 U12 ( .A(b[10]), .Y(n20) );
  XNOR2X1 U13 ( .A(P1[11]), .B(n74), .Y(n128) );
  XNOR2X4 U14 ( .A(b_1), .B(n74), .Y(n57) );
  INVX4 U15 ( .A(b[7]), .Y(n74) );
  INVX1 U16 ( .A(b_2), .Y(n1) );
  BUFX3 U17 ( .A(b[6]), .Y(P1[11]) );
  BUFX3 U18 ( .A(P1[5]), .Y(P2[10]) );
  BUFX8 U19 ( .A(b[8]), .Y(P1[0]) );
  XOR2X2 U20 ( .A(b_0), .B(n9), .Y(n15) );
  INVX1 U21 ( .A(P1[12]), .Y(n8) );
  XNOR2X1 U22 ( .A(n8), .B(P1[3]), .Y(P2[8]) );
  INVX1 U23 ( .A(n15), .Y(n127) );
  XNOR2X1 U24 ( .A(n76), .B(n57), .Y(n59) );
  INVX1 U25 ( .A(b_3), .Y(n30) );
  XOR2X1 U26 ( .A(P2[2]), .B(n59), .Y(n45) );
  XNOR2X1 U27 ( .A(b_0), .B(n16), .Y(n46) );
  XNOR2X1 U28 ( .A(n22), .B(n127), .Y(n114) );
  XNOR2X1 U29 ( .A(n28), .B(b_2), .Y(n98) );
  CLKINVX3 U30 ( .A(b[6]), .Y(n76) );
  INVX1 U31 ( .A(b[9]), .Y(n10) );
  XNOR2X1 U32 ( .A(n37), .B(n66), .Y(P7[8]) );
  XOR2X1 U33 ( .A(n33), .B(n96), .Y(P4[6]) );
  INVX1 U34 ( .A(n3), .Y(n4) );
  XOR2X1 U35 ( .A(P13[1]), .B(n53), .Y(P7[12]) );
  XNOR2X1 U36 ( .A(n1), .B(n104), .Y(P15[4]) );
  XOR2X1 U37 ( .A(n43), .B(n44), .Y(P7[4]) );
  BUFX3 U38 ( .A(P2[8]), .Y(P3[0]) );
  XOR2XL U39 ( .A(n4), .B(n20), .Y(n70) );
  INVX1 U40 ( .A(n74), .Y(P1[12]) );
  INVX1 U41 ( .A(b[10]), .Y(n6) );
  INVX1 U42 ( .A(b_0), .Y(n3) );
  XOR2X1 U43 ( .A(b[12]), .B(n73), .Y(P3[3]) );
  XNOR2X2 U44 ( .A(P1[0]), .B(n76), .Y(n115) );
  XNOR2X2 U45 ( .A(n48), .B(n46), .Y(n97) );
  XNOR2X2 U46 ( .A(b[11]), .B(n26), .Y(n105) );
  XOR2X2 U47 ( .A(n125), .B(n97), .Y(n26) );
  CLKINVX2 U48 ( .A(P1[0]), .Y(n83) );
  XOR2X1 U49 ( .A(b[4]), .B(b[10]), .Y(n33) );
  XOR2X1 U50 ( .A(n36), .B(n51), .Y(P6[8]) );
  XNOR2XL U51 ( .A(b[11]), .B(n36), .Y(P8[3]) );
  XNOR2XL U52 ( .A(n91), .B(P1[0]), .Y(n122) );
  INVX2 U53 ( .A(P1[10]), .Y(n91) );
  BUFX2 U54 ( .A(P16[12]), .Y(P15[7]) );
  XNOR2XL U55 ( .A(n16), .B(b[10]), .Y(n42) );
  XNOR2X1 U56 ( .A(n1), .B(n112), .Y(n95) );
  XNOR2XL U57 ( .A(n1), .B(P1[11]), .Y(n12) );
  XOR2XL U58 ( .A(n1), .B(P1[10]), .Y(n66) );
  XOR2XL U59 ( .A(P1[11]), .B(b[10]), .Y(n107) );
  XNOR2X1 U60 ( .A(P1[11]), .B(n22), .Y(n96) );
  INVX1 U61 ( .A(b[11]), .Y(n2) );
  XNOR2XL U62 ( .A(n2), .B(b[7]), .Y(n117) );
  XNOR2X1 U63 ( .A(b[4]), .B(n2), .Y(n40) );
  INVX1 U64 ( .A(b[11]), .Y(n18) );
  INVX1 U65 ( .A(b[12]), .Y(n5) );
  XNOR2XL U66 ( .A(n22), .B(b[7]), .Y(n68) );
  XNOR2XL U67 ( .A(n22), .B(b_3), .Y(P2[0]) );
  INVX4 U68 ( .A(b[12]), .Y(n22) );
  XOR2X1 U69 ( .A(n20), .B(P1[0]), .Y(n82) );
  XNOR2XL U70 ( .A(n6), .B(b_3), .Y(n61) );
  XNOR2XL U71 ( .A(n20), .B(b[9]), .Y(P1[2]) );
  XNOR2XL U72 ( .A(P1[0]), .B(n9), .Y(P1[1]) );
  BUFX3 U73 ( .A(n30), .Y(n11) );
  XNOR2X1 U74 ( .A(P1[0]), .B(n211), .Y(n112) );
  BUFX3 U75 ( .A(n30), .Y(n211) );
  XOR2XL U76 ( .A(b[10]), .B(n114), .Y(P1[5]) );
  XOR2X1 U77 ( .A(P1[1]), .B(n45), .Y(n43) );
  XNOR2X1 U78 ( .A(n4), .B(n8), .Y(n78) );
  XNOR2XL U79 ( .A(n93), .B(n34), .Y(P9[1]) );
  BUFX3 U80 ( .A(P8[12]), .Y(P7[7]) );
  XNOR2X1 U81 ( .A(n91), .B(P1[11]), .Y(n90) );
  XNOR2X1 U82 ( .A(n93), .B(n65), .Y(P2[11]) );
  XNOR2XL U83 ( .A(n76), .B(n54), .Y(P15[3]) );
  XNOR2XL U84 ( .A(n38), .B(n59), .Y(n100) );
  XNOR2XL U85 ( .A(n62), .B(n97), .Y(n32) );
  XNOR2X1 U86 ( .A(n83), .B(n79), .Y(P11[1]) );
  CLKBUFXL U87 ( .A(P4[6]), .Y(P5[11]) );
  INVXL U88 ( .A(b_1), .Y(n93) );
  XOR2X1 U89 ( .A(P16[4]), .B(P1[1]), .Y(n104) );
  XOR2X1 U90 ( .A(n58), .B(n12), .Y(n85) );
  XOR2XL U91 ( .A(P16[5]), .B(n65), .Y(n102) );
  XOR2XL U92 ( .A(n40), .B(n127), .Y(n88) );
  XOR2X1 U93 ( .A(n4), .B(n55), .Y(P5[3]) );
  XNOR2XL U94 ( .A(n86), .B(n8), .Y(n126) );
  XOR2XL U95 ( .A(n53), .B(n131), .Y(n129) );
  XOR2X1 U96 ( .A(n48), .B(n49), .Y(P7[2]) );
  XOR2X1 U97 ( .A(n42), .B(n43), .Y(P7[5]) );
  XOR2X1 U98 ( .A(n92), .B(n110), .Y(P13[8]) );
  XOR2X1 U99 ( .A(n37), .B(n39), .Y(P8[12]) );
  XOR2X1 U100 ( .A(n55), .B(n56), .Y(P7[10]) );
  XNOR2X1 U101 ( .A(n132), .B(n13), .Y(n116) );
  XNOR2XL U102 ( .A(n18), .B(P1[0]), .Y(n13) );
  XNOR2XL U103 ( .A(n18), .B(b[10]), .Y(n65) );
  XOR2XL U104 ( .A(b[4]), .B(b_3), .Y(P16[4]) );
  INVX1 U105 ( .A(b[4]), .Y(n28) );
  XNOR2XL U106 ( .A(n25), .B(n71), .Y(n24) );
  XNOR2X1 U107 ( .A(P1[10]), .B(b[7]), .Y(n25) );
  XNOR2XL U108 ( .A(b[12]), .B(b_2), .Y(n38) );
  XOR2XL U109 ( .A(n111), .B(n124), .Y(n77) );
  XOR2X1 U110 ( .A(b_1), .B(b[12]), .Y(n111) );
  XNOR2X1 U111 ( .A(P1[5]), .B(b[4]), .Y(n49) );
  XOR2X1 U112 ( .A(n81), .B(n41), .Y(P4[3]) );
  XNOR2XL U113 ( .A(n11), .B(b[9]), .Y(n41) );
  XOR2X1 U114 ( .A(n52), .B(n72), .Y(n55) );
  XOR2X1 U115 ( .A(P6[3]), .B(n29), .Y(P8[7]) );
  XOR2X1 U116 ( .A(P12[3]), .B(n107), .Y(P7[6]) );
  XOR2X1 U117 ( .A(n105), .B(n109), .Y(n54) );
  XOR2XL U118 ( .A(n22), .B(b[10]), .Y(n109) );
  BUFX3 U119 ( .A(P11[6]), .Y(P12[11]) );
  BUFX3 U120 ( .A(P12[12]), .Y(P11[7]) );
  BUFX3 U121 ( .A(P10[0]), .Y(P9[8]) );
  BUFX3 U122 ( .A(P10[5]), .Y(P11[10]) );
  BUFX3 U123 ( .A(P15[6]), .Y(P16[11]) );
  BUFX3 U124 ( .A(P3[5]), .Y(P4[10]) );
  BUFX3 U125 ( .A(P14[11]), .Y(P13[6]) );
  BUFX3 U126 ( .A(P7[4]), .Y(P8[9]) );
  BUFX3 U127 ( .A(P3[6]), .Y(P4[11]) );
  XNOR2X1 U128 ( .A(n83), .B(P9[2]), .Y(P3[5]) );
  XNOR2X1 U129 ( .A(n83), .B(n129), .Y(P12[12]) );
  XNOR2X1 U130 ( .A(n62), .B(P2[5]), .Y(P11[6]) );
  XNOR2X1 U131 ( .A(n76), .B(n102), .Y(P15[6]) );
  XNOR2X1 U132 ( .A(n93), .B(n103), .Y(P14[11]) );
  XOR2X1 U133 ( .A(n119), .B(P2[8]), .Y(P11[9]) );
  XOR2X1 U134 ( .A(n87), .B(n88), .Y(P3[6]) );
  XOR2X1 U135 ( .A(n96), .B(n32), .Y(n31) );
  XNOR2X1 U136 ( .A(n62), .B(n63), .Y(n47) );
  XNOR2X1 U137 ( .A(n91), .B(n92), .Y(P2[3]) );
  XOR2X1 U138 ( .A(n87), .B(n71), .Y(P15[1]) );
  XOR2X1 U139 ( .A(n115), .B(n88), .Y(n69) );
  XOR2X1 U140 ( .A(n118), .B(n119), .Y(n35) );
  XNOR2X1 U141 ( .A(n93), .B(n95), .Y(n14) );
  XNOR2X1 U142 ( .A(n15), .B(n89), .Y(n73) );
  XNOR2X1 U143 ( .A(n83), .B(P2[3]), .Y(P4[2]) );
  XNOR2XL U144 ( .A(n112), .B(n126), .Y(P11[3]) );
  XOR2X1 U145 ( .A(n46), .B(n47), .Y(P7[3]) );
  BUFX3 U146 ( .A(P11[5]), .Y(P12[10]) );
  BUFX3 U147 ( .A(P14[9]), .Y(P13[4]) );
  BUFX3 U148 ( .A(P12[5]), .Y(P13[10]) );
  BUFX3 U149 ( .A(P15[4]), .Y(P16[9]) );
  BUFX3 U150 ( .A(P4[5]), .Y(P5[10]) );
  BUFX3 U151 ( .A(P9[4]), .Y(P10[9]) );
  BUFX3 U152 ( .A(P10[12]), .Y(P9[7]) );
  BUFX3 U153 ( .A(P1[7]), .Y(P2[12]) );
  BUFX3 U154 ( .A(P2[5]), .Y(P3[10]) );
  BUFX3 U155 ( .A(P15[8]), .Y(P16[0]) );
  BUFX3 U156 ( .A(P7[5]), .Y(P8[10]) );
  BUFX3 U157 ( .A(P9[5]), .Y(P10[10]) );
  BUFX3 U158 ( .A(P9[6]), .Y(P10[11]) );
  BUFX3 U159 ( .A(P15[10]), .Y(P14[5]) );
  BUFX3 U160 ( .A(P13[7]), .Y(P14[12]) );
  BUFX3 U161 ( .A(P6[6]), .Y(P7[11]) );
  BUFX3 U162 ( .A(P8[6]), .Y(P9[11]) );
  BUFX3 U163 ( .A(P3[8]), .Y(P4[0]) );
  BUFX3 U164 ( .A(P13[11]), .Y(P12[6]) );
  BUFX3 U165 ( .A(P6[4]), .Y(P7[9]) );
  BUFX3 U166 ( .A(P7[10]), .Y(P6[5]) );
  BUFX3 U167 ( .A(P7[12]), .Y(P6[7]) );
  BUFX3 U168 ( .A(P13[8]), .Y(P14[0]) );
  BUFX3 U169 ( .A(P6[12]), .Y(P5[7]) );
  BUFX3 U170 ( .A(P13[5]), .Y(P14[10]) );
  XOR2X1 U171 ( .A(n90), .B(P1[1]), .Y(P3[11]) );
  XOR2X1 U172 ( .A(P2[2]), .B(n125), .Y(P2[5]) );
  BUFX3 U173 ( .A(P3[11]), .Y(P2[6]) );
  BUFX3 U174 ( .A(P16[10]), .Y(P15[5]) );
  XOR2X1 U175 ( .A(n128), .B(P1[2]), .Y(P3[12]) );
  XNOR2X1 U176 ( .A(n22), .B(n45), .Y(P6[3]) );
  XNOR2X1 U177 ( .A(n83), .B(n65), .Y(P1[3]) );
  XNOR2X1 U178 ( .A(n11), .B(n103), .Y(P16[10]) );
  XOR2X1 U179 ( .A(n4), .B(n121), .Y(P9[2]) );
  XOR2X1 U180 ( .A(n4), .B(P2[2]), .Y(P16[5]) );
  XOR2X1 U181 ( .A(n42), .B(n80), .Y(P5[9]) );
  XOR2X1 U182 ( .A(n42), .B(n99), .Y(P11[11]) );
  XOR2X1 U183 ( .A(b_1), .B(n21), .Y(P16[6]) );
  XOR2X1 U184 ( .A(n58), .B(n78), .Y(P4[7]) );
  XOR2X1 U185 ( .A(n68), .B(n69), .Y(P6[10]) );
  XOR2X1 U186 ( .A(n34), .B(n35), .Y(P9[9]) );
  XNOR2XL U187 ( .A(n6), .B(n21), .Y(P9[5]) );
  XNOR2X1 U188 ( .A(n20), .B(n85), .Y(P13[7]) );
  XNOR2X1 U189 ( .A(n6), .B(n104), .Y(P15[10]) );
  XNOR2X1 U190 ( .A(n2), .B(n100), .Y(P15[0]) );
  XNOR2X1 U191 ( .A(n2), .B(n19), .Y(P9[6]) );
  XNOR2X1 U192 ( .A(n28), .B(n54), .Y(P6[6]) );
  XNOR2X1 U193 ( .A(n28), .B(n17), .Y(P13[9]) );
  XNOR2X1 U194 ( .A(n28), .B(n31), .Y(P8[6]) );
  XNOR2X1 U195 ( .A(n76), .B(n77), .Y(P5[0]) );
  XNOR2X1 U196 ( .A(n11), .B(n80), .Y(P10[8]) );
  XNOR2X1 U197 ( .A(n11), .B(P3[12]), .Y(P11[8]) );
  XNOR2XL U198 ( .A(n11), .B(n129), .Y(P12[9]) );
  XNOR2X1 U199 ( .A(n10), .B(n67), .Y(P6[11]) );
  XNOR2X1 U200 ( .A(n8), .B(P9[1]), .Y(P3[4]) );
  XNOR2X1 U201 ( .A(n11), .B(n85), .Y(P3[8]) );
  XNOR2X1 U202 ( .A(n10), .B(n94), .Y(P1[4]) );
  XNOR2X1 U203 ( .A(n10), .B(n108), .Y(P14[4]) );
  XNOR2X1 U204 ( .A(n10), .B(n102), .Y(P14[6]) );
  XOR2XL U205 ( .A(n98), .B(n116), .Y(P12[8]) );
  XOR2X1 U206 ( .A(n61), .B(n47), .Y(P5[8]) );
  XOR2X1 U207 ( .A(P9[1]), .B(n122), .Y(P12[5]) );
  XOR2X1 U208 ( .A(P9[2]), .B(n120), .Y(P13[11]) );
  XNOR2XL U209 ( .A(n10), .B(P1[11]), .Y(n120) );
  XOR2X1 U210 ( .A(n35), .B(n117), .Y(P13[12]) );
  XOR2X1 U211 ( .A(n121), .B(n117), .Y(P11[12]) );
  XOR2X1 U212 ( .A(P10[3]), .B(n58), .Y(P6[4]) );
  XNOR2X1 U213 ( .A(P8[1]), .B(n70), .Y(P11[5]) );
  XOR2X1 U214 ( .A(n24), .B(n61), .Y(P5[4]) );
  XOR2X1 U215 ( .A(n64), .B(n65), .Y(P6[12]) );
  XOR2X1 U216 ( .A(n4), .B(n104), .Y(P13[5]) );
  XNOR2X1 U217 ( .A(n18), .B(n78), .Y(n110) );
  XNOR2XL U218 ( .A(n211), .B(P1[11]), .Y(n39) );
  XOR2X1 U219 ( .A(n26), .B(n27), .Y(P8[8]) );
  XOR2XL U220 ( .A(n53), .B(n89), .Y(n67) );
  XNOR2X1 U221 ( .A(n83), .B(n50), .Y(n94) );
  XNOR2X1 U222 ( .A(n6), .B(P14[2]), .Y(P13[2]) );
  XNOR2X1 U223 ( .A(n76), .B(n34), .Y(n131) );
  XNOR2X1 U224 ( .A(n2), .B(n115), .Y(n71) );
  XNOR2X1 U225 ( .A(n28), .B(n94), .Y(n80) );
  XNOR2X1 U226 ( .A(n6), .B(n23), .Y(n103) );
  XNOR2X1 U227 ( .A(n8), .B(n98), .Y(n84) );
  XNOR2X1 U228 ( .A(n10), .B(n58), .Y(P10[2]) );
  XNOR2X1 U229 ( .A(n10), .B(n68), .Y(n63) );
  XOR2X1 U230 ( .A(b_0), .B(n90), .Y(n21) );
  XNOR2X1 U231 ( .A(n57), .B(n82), .Y(n89) );
  XOR2X1 U232 ( .A(P16[4]), .B(n128), .Y(P8[1]) );
  XNOR2X1 U233 ( .A(n93), .B(n18), .Y(n62) );
  XNOR2X1 U234 ( .A(n6), .B(n84), .Y(P16[2]) );
  XNOR2X1 U235 ( .A(n11), .B(n99), .Y(P16[1]) );
  XNOR2X1 U236 ( .A(n8), .B(n14), .Y(P16[8]) );
  XNOR2X1 U237 ( .A(n76), .B(P2[0]), .Y(n92) );
  XNOR2X1 U238 ( .A(n211), .B(n42), .Y(n121) );
  XNOR2XL U239 ( .A(n28), .B(b_0), .Y(n119) );
  XNOR2X1 U240 ( .A(P1[0]), .B(n74), .Y(n125) );
  XNOR2X1 U241 ( .A(P14[1]), .B(n10), .Y(P13[1]) );
  XNOR2X1 U242 ( .A(b_0), .B(n83), .Y(n124) );
  XOR2X1 U243 ( .A(b_1), .B(n61), .Y(n118) );
  XOR2X1 U244 ( .A(n75), .B(n118), .Y(P10[3]) );
  XOR2X1 U245 ( .A(n105), .B(n10), .Y(P12[3]) );
  XNOR2X1 U246 ( .A(n83), .B(n100), .Y(P15[8]) );
  XNOR2X1 U247 ( .A(P16[6]), .B(n50), .Y(n101) );
  XNOR2X1 U248 ( .A(n9), .B(P2[2]), .Y(n23) );
  XNOR2X1 U249 ( .A(n8), .B(n95), .Y(n108) );
  XNOR2X1 U250 ( .A(n211), .B(P10[2]), .Y(n79) );
  XNOR2X1 U251 ( .A(n8), .B(n77), .Y(n17) );
  XNOR2X1 U252 ( .A(b_1), .B(n211), .Y(n87) );
  XOR2X1 U253 ( .A(n4), .B(n59), .Y(n19) );
  XNOR2X1 U254 ( .A(b_1), .B(n53), .Y(n132) );
  XOR2X1 U255 ( .A(n52), .B(n44), .Y(P13[3]) );
  BUFX3 U256 ( .A(P3[9]), .Y(P2[4]) );
  XOR2X1 U257 ( .A(n4), .B(P1[3]), .Y(P3[2]) );
  XOR2X1 U258 ( .A(n4), .B(P2[5]), .Y(P8[2]) );
  XNOR2X1 U259 ( .A(n24), .B(n106), .Y(P9[3]) );
  XOR2X1 U260 ( .A(n1), .B(b_1), .Y(n106) );
  BUFX3 U261 ( .A(P2[11]), .Y(P1[6]) );
  XNOR2X1 U262 ( .A(n8), .B(n31), .Y(P16[3]) );
  XOR2X1 U263 ( .A(n58), .B(n84), .Y(n81) );
  XOR2XL U264 ( .A(n132), .B(n33), .Y(n86) );
  XNOR2X1 U265 ( .A(P1[11]), .B(n49), .Y(P11[2]) );
  BUFX3 U266 ( .A(P4[7]), .Y(P5[12]) );
  XOR2X1 U267 ( .A(P15[4]), .B(n60), .Y(P6[2]) );
  BUFX3 U268 ( .A(P13[9]), .Y(P12[4]) );
  BUFX3 U269 ( .A(P10[8]), .Y(P11[0]) );
  BUFX3 U270 ( .A(P13[12]), .Y(P12[7]) );
  BUFX3 U271 ( .A(P8[5]), .Y(P9[10]) );
  XNOR2X1 U272 ( .A(n11), .B(n69), .Y(P12[1]) );
  BUFX3 U273 ( .A(P11[9]), .Y(P10[4]) );
  BUFX3 U274 ( .A(P11[12]), .Y(P10[7]) );
  BUFX3 U275 ( .A(P8[8]), .Y(P9[0]) );
  BUFX3 U276 ( .A(P5[8]), .Y(P6[0]) );
  BUFX3 U277 ( .A(P5[4]), .Y(P6[9]) );
  BUFX3 U278 ( .A(P6[10]), .Y(P5[5]) );
  BUFX3 U279 ( .A(P5[0]), .Y(P4[8]) );
  BUFX3 U280 ( .A(P3[12]), .Y(P2[7]) );
  BUFX3 U281 ( .A(P14[4]), .Y(P15[9]) );
  BUFX3 U282 ( .A(P6[8]), .Y(P7[0]) );
  BUFX3 U283 ( .A(P11[11]), .Y(P10[6]) );
  BUFX3 U284 ( .A(P6[11]), .Y(P5[6]) );
  BUFX3 U285 ( .A(P5[9]), .Y(P4[4]) );
  BUFX3 U286 ( .A(P7[8]), .Y(P8[0]) );
  XNOR2X1 U287 ( .A(n2), .B(n67), .Y(P14[3]) );
  BUFX3 U288 ( .A(P11[8]), .Y(P12[0]) );
  BUFX3 U289 ( .A(P12[9]), .Y(P11[4]) );
  BUFX3 U290 ( .A(P9[9]), .Y(P8[4]) );
  XOR2X1 U291 ( .A(P15[4]), .B(n50), .Y(P7[1]) );
  BUFX3 U292 ( .A(P3[4]), .Y(P4[9]) );
  XNOR2X1 U293 ( .A(n6), .B(n63), .Y(P3[1]) );
  XNOR2X1 U294 ( .A(n28), .B(P2[0]), .Y(P2[1]) );
  BUFX3 U295 ( .A(P1[4]), .Y(P2[9]) );
  BUFX3 U296 ( .A(P15[0]), .Y(P14[8]) );
  BUFX3 U297 ( .A(P14[6]), .Y(P15[11]) );
  BUFX3 U298 ( .A(P12[8]), .Y(P13[0]) );
  BUFX3 U299 ( .A(P2[0]), .Y(P1[8]) );
  BUFX3 U300 ( .A(P3[7]), .Y(P4[12]) );
  BUFX3 U301 ( .A(P15[12]), .Y(P14[7]) );
  BUFX3 U302 ( .A(P7[6]), .Y(P8[11]) );
  BUFX3 U303 ( .A(P8[7]), .Y(P9[12]) );
  XNOR2X1 U304 ( .A(n4), .B(n211), .Y(n44) );
  XNOR2XL U305 ( .A(n6), .B(P1[10]), .Y(n60) );
  XOR2X1 U306 ( .A(P1[10]), .B(b[11]), .Y(n58) );
  XOR2X1 U307 ( .A(P1[10]), .B(b[4]), .Y(P2[2]) );
  XOR2X1 U308 ( .A(b_2), .B(P4[6]), .Y(n52) );
  XNOR2X1 U309 ( .A(b[10]), .B(n101), .Y(P15[12]) );
  XNOR2XL U310 ( .A(n133), .B(n96), .Y(n99) );
  XOR2X1 U311 ( .A(b[4]), .B(P15[1]), .Y(P14[1]) );
  XNOR2X1 U312 ( .A(P1[10]), .B(b_3), .Y(n48) );
  XOR2X1 U313 ( .A(b[12]), .B(n64), .Y(n75) );
  XOR2X1 U314 ( .A(n113), .B(n98), .Y(P15[2]) );
  XOR2X1 U315 ( .A(b[7]), .B(n114), .Y(n113) );
  CLKBUFXL U316 ( .A(b[4]), .Y(P1[9]) );
  XNOR2X1 U317 ( .A(n10), .B(b[11]), .Y(n72) );
  XNOR2X1 U318 ( .A(n22), .B(n108), .Y(P14[9]) );
  XNOR2X1 U319 ( .A(n22), .B(P8[1]), .Y(P3[9]) );
  XNOR2X1 U320 ( .A(n22), .B(n79), .Y(P4[5]) );
  XNOR2X1 U321 ( .A(n5), .B(n81), .Y(P4[1]) );
  XNOR2X1 U322 ( .A(n22), .B(n23), .Y(P9[4]) );
  XNOR2X1 U323 ( .A(n18), .B(b[12]), .Y(n50) );
  XNOR2X1 U324 ( .A(P15[2]), .B(n91), .Y(P14[2]) );
  XNOR2XL U325 ( .A(n8), .B(n75), .Y(P5[1]) );
  XNOR2X1 U326 ( .A(n1), .B(n19), .Y(P16[7]) );
  XNOR2X1 U327 ( .A(n1), .B(n50), .Y(P1[7]) );
  XNOR2X1 U328 ( .A(b_2), .B(n86), .Y(P3[7]) );
  XNOR2X1 U329 ( .A(n1), .B(n17), .Y(P10[12]) );
  XNOR2X1 U330 ( .A(n11), .B(b_2), .Y(n29) );
  XNOR2XL U331 ( .A(n14), .B(n15), .Y(P10[0]) );
  XNOR2X1 U332 ( .A(n15), .B(n116), .Y(P10[5]) );
  XNOR2X1 U333 ( .A(b[9]), .B(n126), .Y(P12[2]) );
  XNOR2X1 U334 ( .A(P1[10]), .B(b[9]), .Y(n51) );
  XNOR2XL U335 ( .A(b_1), .B(b[9]), .Y(n133) );
  XNOR2XL U336 ( .A(n11), .B(n73), .Y(P5[2]) );
  XOR2X1 U337 ( .A(n57), .B(P15[4]), .Y(P6[1]) );
  XNOR2X1 U338 ( .A(b[7]), .B(n101), .Y(P16[12]) );
  XNOR2XL U339 ( .A(n211), .B(n57), .Y(n56) );
endmodule


module multiplier_column4_p16 ( b, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, 
        P11, P12, P13, P14, P15, P16 );
  input [12:0] b;
  output [12:0] P1;
  output [12:0] P2;
  output [12:0] P3;
  output [12:0] P4;
  output [12:0] P5;
  output [12:0] P6;
  output [12:0] P7;
  output [12:0] P8;
  output [12:0] P9;
  output [12:0] P10;
  output [12:0] P11;
  output [12:0] P12;
  output [12:0] P13;
  output [12:0] P14;
  output [12:0] P15;
  output [12:0] P16;
  wire   b_12, b_11, b_10, n240, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n48, n49, n50, n51, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n86, n87, n88, n89, n90, n91, n92, n95, n96, n97, n101, n102,
         n103, n104, n106, n107, n108, n110, n111, n112, n114, n117, n118,
         n119, n120, n122, n123, n1, n2, n3, n5, n6, n7, n8, n9, n10, n12, n13,
         n14, n47, n52, n69, n85, n93, n94, n98, n99, n100, n105, n109, n113,
         n116, n121, n124, n125, n126, n127, n128, n129, n130, n131, n222,
         n223;
  assign b_12 = b[12];
  assign b_11 = b[11];
  assign b_10 = b[10];

  INVX1 U1 ( .A(n8), .Y(n1) );
  INVX2 U2 ( .A(b[2]), .Y(n26) );
  DLY1X1 U3 ( .A(P5[4]), .Y(P7[12]) );
  DLY1X1 U4 ( .A(P5[4]), .Y(P6[8]) );
  NAND2X4 U5 ( .A(b_10), .B(n26), .Y(n9) );
  INVX1 U6 ( .A(b_12), .Y(n2) );
  BUFX3 U7 ( .A(b[0]), .Y(n222) );
  XOR2X1 U8 ( .A(n48), .B(n49), .Y(n240) );
  OAI2BB1X2 U9 ( .A0N(n240), .A1N(n85), .B0(n93), .Y(n27) );
  OAI2BB1X2 U10 ( .A0N(n67), .A1N(n40), .B0(n52), .Y(P1[3]) );
  XOR2X1 U11 ( .A(n28), .B(n31), .Y(P9[9]) );
  OAI2BB1X1 U12 ( .A0N(n30), .A1N(P2[2]), .B0(n99), .Y(n119) );
  NAND2BX1 U13 ( .AN(n102), .B(P3[11]), .Y(n13) );
  OAI2BB1X2 U14 ( .A0N(n126), .A1N(n5), .B0(n7), .Y(P8[12]) );
  INVXL U15 ( .A(P4[3]), .Y(n5) );
  XOR2X2 U16 ( .A(P1[12]), .B(P2[1]), .Y(n64) );
  OAI2BB1X2 U17 ( .A0N(n35), .A1N(P1[2]), .B0(n94), .Y(P1[5]) );
  XOR2X1 U18 ( .A(n50), .B(n19), .Y(P4[3]) );
  NAND2X1 U19 ( .A(n13), .B(n14), .Y(P14[11]) );
  XNOR2X4 U20 ( .A(n2), .B(n32), .Y(n112) );
  NAND2X4 U21 ( .A(n9), .B(n10), .Y(n32) );
  NAND2X2 U22 ( .A(n8), .B(b[2]), .Y(n10) );
  XNOR2XL U23 ( .A(P1[11]), .B(n37), .Y(P8[1]) );
  INVX8 U24 ( .A(P1[12]), .Y(n68) );
  XNOR2X4 U25 ( .A(n67), .B(b_11), .Y(n90) );
  INVX4 U26 ( .A(b[9]), .Y(n67) );
  XNOR2X2 U27 ( .A(b_10), .B(n56), .Y(P1[2]) );
  XOR2X2 U28 ( .A(b[9]), .B(n64), .Y(P2[4]) );
  INVX1 U29 ( .A(n240), .Y(n69) );
  XNOR2X1 U30 ( .A(P4[1]), .B(n222), .Y(n50) );
  INVX1 U31 ( .A(b_12), .Y(n55) );
  CLKINVX3 U32 ( .A(b[3]), .Y(n30) );
  BUFX3 U33 ( .A(P1[5]), .Y(P2[9]) );
  CLKBUFX8 U34 ( .A(b[6]), .Y(P1[10]) );
  BUFX4 U35 ( .A(b[5]), .Y(P2[0]) );
  XOR2X1 U36 ( .A(P1[5]), .B(P2[11]), .Y(n48) );
  XNOR2X2 U37 ( .A(n65), .B(P1[10]), .Y(P2[1]) );
  BUFX3 U38 ( .A(P1[5]), .Y(P3[0]) );
  XOR2X2 U39 ( .A(P2[12]), .B(n119), .Y(P10[1]) );
  XNOR2X2 U40 ( .A(n120), .B(n56), .Y(P11[2]) );
  XOR2X2 U41 ( .A(P1[12]), .B(P1[3]), .Y(P3[11]) );
  XNOR2X1 U42 ( .A(n8), .B(P1[10]), .Y(n16) );
  XNOR2X1 U43 ( .A(n1), .B(P1[11]), .Y(n82) );
  CLKBUFX8 U44 ( .A(b[7]), .Y(P1[11]) );
  XNOR2X4 U45 ( .A(n223), .B(n112), .Y(n81) );
  XOR2X1 U46 ( .A(n63), .B(n22), .Y(P15[3]) );
  XOR2X1 U47 ( .A(n28), .B(n29), .Y(P9[10]) );
  XNOR2X1 U48 ( .A(n30), .B(n96), .Y(P16[0]) );
  BUFX3 U49 ( .A(P15[10]), .Y(P14[6]) );
  INVX1 U50 ( .A(P2[2]), .Y(n98) );
  BUFX3 U51 ( .A(b[2]), .Y(n3) );
  XNOR2X1 U52 ( .A(n74), .B(n91), .Y(n102) );
  XOR2X1 U53 ( .A(P13[7]), .B(n32), .Y(n28) );
  NAND2X1 U54 ( .A(P1[0]), .B(n47), .Y(n52) );
  INVX4 U55 ( .A(P2[0]), .Y(n65) );
  INVXL U56 ( .A(n69), .Y(P6[7]) );
  XNOR2X1 U57 ( .A(n68), .B(n96), .Y(P13[4]) );
  INVX4 U58 ( .A(b_10), .Y(n8) );
  INVX4 U59 ( .A(b[1]), .Y(n35) );
  INVX1 U60 ( .A(n67), .Y(P1[0]) );
  XNOR2X1 U61 ( .A(n81), .B(n65), .Y(n34) );
  XNOR2X1 U62 ( .A(n19), .B(P1[12]), .Y(n104) );
  XOR2X4 U63 ( .A(P5[4]), .B(n62), .Y(P12[3]) );
  XNOR2X2 U64 ( .A(n65), .B(b[3]), .Y(n62) );
  INVX4 U65 ( .A(P1[10]), .Y(n42) );
  BUFX3 U66 ( .A(P4[7]), .Y(P5[11]) );
  XNOR2X1 U67 ( .A(n26), .B(n40), .Y(P2[10]) );
  INVX1 U68 ( .A(n40), .Y(n47) );
  XNOR2X2 U69 ( .A(n56), .B(b_12), .Y(n40) );
  XOR2X1 U70 ( .A(P2[10]), .B(n108), .Y(P13[1]) );
  XOR2X2 U71 ( .A(n21), .B(P12[3]), .Y(P9[12]) );
  XOR2X2 U72 ( .A(P1[11]), .B(n222), .Y(n21) );
  XNOR2XL U73 ( .A(n67), .B(n32), .Y(n123) );
  XNOR2X1 U74 ( .A(n32), .B(n50), .Y(P7[10]) );
  XNOR2X1 U75 ( .A(n30), .B(b_12), .Y(P2[11]) );
  XOR2X2 U76 ( .A(n22), .B(n27), .Y(P10[12]) );
  XNOR2X1 U77 ( .A(P1[11]), .B(n101), .Y(P14[1]) );
  XNOR2XL U78 ( .A(n3), .B(P1[11]), .Y(n88) );
  XNOR2XL U79 ( .A(n67), .B(P1[11]), .Y(n49) );
  XNOR2X4 U80 ( .A(n42), .B(P1[11]), .Y(P2[2]) );
  BUFX3 U81 ( .A(b[4]), .Y(P2[12]) );
  BUFX3 U82 ( .A(b[4]), .Y(n223) );
  NAND2XL U83 ( .A(P4[3]), .B(n6), .Y(n7) );
  INVXL U84 ( .A(n126), .Y(n6) );
  BUFX2 U85 ( .A(P8[12]), .Y(P7[8]) );
  BUFX2 U86 ( .A(P8[12]), .Y(P6[4]) );
  XOR2XL U87 ( .A(P4[10]), .B(n90), .Y(n131) );
  XNOR2X4 U88 ( .A(n68), .B(n90), .Y(n71) );
  XOR2X1 U89 ( .A(n62), .B(n90), .Y(n89) );
  XOR2X4 U90 ( .A(n101), .B(n56), .Y(P5[4]) );
  INVX2 U91 ( .A(P1[2]), .Y(n73) );
  NAND2X2 U92 ( .A(n12), .B(n102), .Y(n14) );
  NAND2X2 U93 ( .A(n13), .B(n14), .Y(P13[7]) );
  CLKINVX3 U94 ( .A(P3[11]), .Y(n12) );
  XOR2XL U95 ( .A(n62), .B(P1[3]), .Y(P5[5]) );
  NAND2X1 U96 ( .A(b[1]), .B(n73), .Y(n94) );
  NAND2X1 U97 ( .A(n69), .B(n33), .Y(n93) );
  INVX1 U98 ( .A(n33), .Y(n85) );
  XOR2XL U99 ( .A(n20), .B(n21), .Y(P9[5]) );
  NAND2X1 U100 ( .A(b[3]), .B(n98), .Y(n99) );
  XOR2X1 U101 ( .A(P15[3]), .B(n16), .Y(P10[11]) );
  XNOR2XL U102 ( .A(n42), .B(n222), .Y(n107) );
  XNOR2X1 U103 ( .A(n42), .B(P2[12]), .Y(n33) );
  BUFX3 U104 ( .A(P9[4]), .Y(P10[8]) );
  CLKBUFXL U105 ( .A(P3[7]), .Y(P4[11]) );
  CLKBUFXL U106 ( .A(P9[12]), .Y(P8[8]) );
  XNOR2X1 U107 ( .A(P4[2]), .B(n91), .Y(n51) );
  XNOR2X4 U108 ( .A(n81), .B(n68), .Y(n101) );
  XNOR2X1 U109 ( .A(n74), .B(P1[12]), .Y(n22) );
  XOR2X1 U110 ( .A(P1[1]), .B(P2[2]), .Y(P2[5]) );
  XNOR2X1 U111 ( .A(n19), .B(P2[12]), .Y(n31) );
  XNOR2X1 U112 ( .A(n35), .B(P1[10]), .Y(n109) );
  XOR2X1 U113 ( .A(n95), .B(n125), .Y(n23) );
  XOR2X1 U114 ( .A(n26), .B(P2[0]), .Y(n125) );
  XNOR2X1 U115 ( .A(b[9]), .B(n42), .Y(n83) );
  XOR2XL U116 ( .A(P2[0]), .B(b_11), .Y(n128) );
  XNOR2X1 U117 ( .A(b[9]), .B(b[3]), .Y(n124) );
  CLKBUFXL U118 ( .A(P9[5]), .Y(P11[0]) );
  CLKBUFXL U119 ( .A(P9[5]), .Y(P10[9]) );
  CLKBUFXL U120 ( .A(P10[12]), .Y(P8[4]) );
  INVXL U121 ( .A(P10[1]), .Y(n95) );
  XNOR2XL U122 ( .A(n19), .B(P2[1]), .Y(n18) );
  XOR2X1 U123 ( .A(n22), .B(n23), .Y(P9[4]) );
  CLKBUFXL U124 ( .A(P4[10]), .Y(P3[6]) );
  CLKBUFXL U125 ( .A(P6[12]), .Y(P5[8]) );
  CLKBUFXL U126 ( .A(P3[11]), .Y(P2[7]) );
  CLKINVX3 U127 ( .A(n223), .Y(n61) );
  XOR2X1 U128 ( .A(n92), .B(n100), .Y(P13[10]) );
  XNOR2XL U129 ( .A(n55), .B(P1[12]), .Y(n100) );
  XOR2X1 U130 ( .A(n24), .B(n105), .Y(P6[0]) );
  XNOR2XL U131 ( .A(n35), .B(P1[11]), .Y(n105) );
  XOR2X1 U132 ( .A(P12[2]), .B(n109), .Y(P13[0]) );
  XNOR2X1 U133 ( .A(n114), .B(n113), .Y(n87) );
  XOR2X1 U134 ( .A(n74), .B(n104), .Y(n113) );
  XOR2XL U135 ( .A(n77), .B(P2[1]), .Y(n72) );
  XOR2X1 U136 ( .A(n97), .B(n116), .Y(P14[4]) );
  XNOR2XL U137 ( .A(n61), .B(P1[12]), .Y(n116) );
  XNOR2XL U138 ( .A(n30), .B(P2[1]), .Y(n38) );
  XNOR2XL U139 ( .A(n74), .B(P2[12]), .Y(n103) );
  XNOR2X1 U140 ( .A(n84), .B(n121), .Y(P15[5]) );
  XOR2X1 U141 ( .A(n68), .B(n86), .Y(n121) );
  XNOR2XL U142 ( .A(n30), .B(P1[10]), .Y(n29) );
  CLKBUFXL U143 ( .A(P2[4]), .Y(P4[12]) );
  XOR2X1 U144 ( .A(n23), .B(n114), .Y(P11[11]) );
  CLKBUFXL U145 ( .A(P2[4]), .Y(P3[8]) );
  CLKBUFXL U146 ( .A(P2[12]), .Y(P1[8]) );
  XNOR2XL U147 ( .A(n118), .B(n119), .Y(n76) );
  XOR2X1 U148 ( .A(n127), .B(n106), .Y(n96) );
  XNOR2X1 U149 ( .A(n124), .B(n22), .Y(n79) );
  CLKBUFXL U150 ( .A(P6[7]), .Y(P7[11]) );
  BUFX3 U151 ( .A(P11[4]), .Y(P12[8]) );
  BUFX3 U152 ( .A(P3[12]), .Y(P2[8]) );
  BUFX3 U153 ( .A(P3[12]), .Y(P1[4]) );
  BUFX3 U154 ( .A(P11[4]), .Y(P13[12]) );
  BUFX3 U155 ( .A(P9[4]), .Y(P11[12]) );
  CLKBUFXL U156 ( .A(P10[12]), .Y(P9[8]) );
  BUFX3 U157 ( .A(P16[8]), .Y(P15[4]) );
  BUFX3 U158 ( .A(P13[11]), .Y(P12[7]) );
  BUFX3 U159 ( .A(P10[11]), .Y(P9[7]) );
  BUFX3 U160 ( .A(P3[10]), .Y(P2[6]) );
  XNOR2X1 U161 ( .A(n42), .B(n117), .Y(P11[4]) );
  XNOR2X1 U162 ( .A(n74), .B(n75), .Y(P3[12]) );
  XNOR2X1 U163 ( .A(n61), .B(P2[3]), .Y(P3[7]) );
  XNOR2X1 U164 ( .A(n73), .B(n104), .Y(P3[10]) );
  XNOR2X1 U165 ( .A(n61), .B(n87), .Y(P16[8]) );
  XNOR2X1 U166 ( .A(n73), .B(n70), .Y(P9[3]) );
  XOR2X1 U167 ( .A(P2[10]), .B(n31), .Y(n66) );
  XNOR2X1 U168 ( .A(n97), .B(n107), .Y(n37) );
  XNOR2X1 U169 ( .A(n61), .B(n106), .Y(P13[11]) );
  XOR2X1 U170 ( .A(n17), .B(n18), .Y(P10[10]) );
  XNOR2X1 U171 ( .A(n25), .B(n60), .Y(n43) );
  XNOR2X1 U172 ( .A(n65), .B(n104), .Y(P2[3]) );
  XNOR2X1 U173 ( .A(n65), .B(n58), .Y(P16[5]) );
  XNOR2X1 U174 ( .A(n25), .B(n107), .Y(n70) );
  XOR2X1 U175 ( .A(n34), .B(n49), .Y(n39) );
  XNOR2X1 U176 ( .A(n74), .B(P3[7]), .Y(P10[2]) );
  BUFX3 U177 ( .A(P14[10]), .Y(P13[6]) );
  BUFX3 U178 ( .A(P12[5]), .Y(P13[9]) );
  BUFX3 U179 ( .A(P15[0]), .Y(P14[9]) );
  BUFX3 U180 ( .A(P16[10]), .Y(P15[6]) );
  BUFX3 U181 ( .A(P10[10]), .Y(P9[6]) );
  BUFX3 U182 ( .A(P2[5]), .Y(P4[0]) );
  XOR2X1 U183 ( .A(n16), .B(n66), .Y(P10[3]) );
  XNOR2X1 U184 ( .A(n25), .B(P12[5]), .Y(P9[1]) );
  XNOR2X1 U185 ( .A(n65), .B(n66), .Y(P5[1]) );
  XNOR2X1 U186 ( .A(n42), .B(n43), .Y(P7[3]) );
  XOR2X1 U187 ( .A(n22), .B(n45), .Y(P15[1]) );
  XOR2X1 U188 ( .A(P9[3]), .B(n31), .Y(P13[3]) );
  BUFX3 U189 ( .A(P8[0]), .Y(P6[5]) );
  BUFX3 U190 ( .A(P8[0]), .Y(P7[9]) );
  BUFX3 U191 ( .A(P12[12]), .Y(P11[8]) );
  BUFX3 U192 ( .A(P12[12]), .Y(P10[4]) );
  BUFX3 U193 ( .A(P14[4]), .Y(P16[12]) );
  BUFX3 U194 ( .A(P15[7]), .Y(P16[11]) );
  BUFX3 U195 ( .A(P15[5]), .Y(P16[9]) );
  BUFX3 U196 ( .A(P2[5]), .Y(P3[9]) );
  BUFX3 U197 ( .A(P12[5]), .Y(P14[0]) );
  BUFX3 U198 ( .A(P16[0]), .Y(P14[5]) );
  BUFX3 U199 ( .A(P16[0]), .Y(P15[9]) );
  BUFX3 U200 ( .A(P13[0]), .Y(P12[9]) );
  BUFX3 U201 ( .A(P13[0]), .Y(P11[5]) );
  BUFX3 U202 ( .A(P14[4]), .Y(P15[8]) );
  BUFX3 U203 ( .A(P13[4]), .Y(P14[8]) );
  BUFX3 U204 ( .A(P13[4]), .Y(P15[12]) );
  BUFX3 U205 ( .A(P5[0]), .Y(P4[9]) );
  BUFX3 U206 ( .A(P5[0]), .Y(P3[5]) );
  BUFX3 U207 ( .A(P11[9]), .Y(P12[0]) );
  BUFX3 U208 ( .A(P11[9]), .Y(P10[5]) );
  BUFX3 U209 ( .A(P15[0]), .Y(P13[5]) );
  BUFX3 U210 ( .A(P12[4]), .Y(P14[12]) );
  BUFX3 U211 ( .A(P12[4]), .Y(P13[8]) );
  BUFX3 U212 ( .A(P13[10]), .Y(P12[6]) );
  BUFX3 U213 ( .A(P10[6]), .Y(P11[10]) );
  BUFX3 U214 ( .A(P15[11]), .Y(P14[7]) );
  BUFX3 U215 ( .A(P12[10]), .Y(P11[6]) );
  BUFX3 U216 ( .A(P11[7]), .Y(P12[11]) );
  BUFX3 U217 ( .A(P11[11]), .Y(P10[7]) );
  CLKBUFXL U218 ( .A(P2[10]), .Y(P1[6]) );
  XNOR2X1 U219 ( .A(n82), .B(P3[2]), .Y(P12[5]) );
  XOR2X1 U220 ( .A(n64), .B(P2[11]), .Y(P5[2]) );
  XNOR2X1 U221 ( .A(n30), .B(n72), .Y(P5[0]) );
  XOR2X1 U222 ( .A(n117), .B(n122), .Y(P11[9]) );
  XNOR2X1 U223 ( .A(n30), .B(P2[5]), .Y(P15[0]) );
  XOR2X1 U224 ( .A(n83), .B(P3[1]), .Y(P12[4]) );
  XOR2X1 U225 ( .A(n83), .B(P11[1]), .Y(P16[10]) );
  XNOR2X1 U226 ( .A(P10[1]), .B(n55), .Y(P4[10]) );
  XOR2X1 U227 ( .A(P1[1]), .B(n78), .Y(n58) );
  XNOR2X1 U228 ( .A(n55), .B(P1[1]), .Y(n75) );
  XNOR2X1 U229 ( .A(n55), .B(n86), .Y(n106) );
  XNOR2X1 U230 ( .A(n30), .B(n49), .Y(n60) );
  XNOR2X1 U231 ( .A(n61), .B(n53), .Y(n41) );
  XOR2X1 U232 ( .A(n59), .B(n111), .Y(P11[1]) );
  XOR2X1 U233 ( .A(P2[4]), .B(n41), .Y(n20) );
  XOR2X1 U234 ( .A(n20), .B(n40), .Y(P9[0]) );
  XNOR2X1 U235 ( .A(n95), .B(n59), .Y(P15[10]) );
  XNOR2X1 U236 ( .A(n110), .B(n37), .Y(P10[6]) );
  XNOR2X1 U237 ( .A(n68), .B(n80), .Y(P15[11]) );
  XNOR2X1 U238 ( .A(n26), .B(n87), .Y(P12[10]) );
  XOR2X1 U239 ( .A(n79), .B(n84), .Y(P11[7]) );
  XNOR2X1 U240 ( .A(n65), .B(n59), .Y(n117) );
  XOR2X1 U241 ( .A(n83), .B(n92), .Y(n45) );
  INVX1 U242 ( .A(b[7]), .Y(n19) );
  XOR2X1 U243 ( .A(P3[10]), .B(n103), .Y(P14[10]) );
  INVX1 U244 ( .A(n222), .Y(n74) );
  XOR2X1 U245 ( .A(n62), .B(P9[3]), .Y(P16[2]) );
  XNOR2X1 U246 ( .A(n30), .B(n80), .Y(P16[3]) );
  XNOR2X1 U247 ( .A(n8), .B(n72), .Y(P16[6]) );
  XNOR2X1 U248 ( .A(n61), .B(n79), .Y(P16[4]) );
  XNOR2X1 U249 ( .A(n222), .B(n39), .Y(P16[1]) );
  XNOR2X1 U250 ( .A(n57), .B(n76), .Y(n36) );
  XOR2X1 U251 ( .A(P1[10]), .B(n71), .Y(P4[1]) );
  XOR2X1 U252 ( .A(P1[11]), .B(n75), .Y(P4[2]) );
  XNOR2X1 U253 ( .A(P1[12]), .B(n51), .Y(P8[0]) );
  XOR2XL U254 ( .A(n62), .B(n71), .Y(P14[2]) );
  XNOR2X1 U255 ( .A(n57), .B(n58), .Y(n17) );
  XNOR2X1 U256 ( .A(n55), .B(n16), .Y(P12[1]) );
  BUFX3 U257 ( .A(P3[4]), .Y(P5[12]) );
  XOR2X1 U258 ( .A(n43), .B(n59), .Y(P6[1]) );
  XNOR2X1 U259 ( .A(n55), .B(n60), .Y(P13[2]) );
  XNOR2XL U260 ( .A(n61), .B(n63), .Y(P5[3]) );
  XNOR2XL U261 ( .A(n61), .B(n48), .Y(P3[3]) );
  XNOR2X1 U262 ( .A(P2[12]), .B(n51), .Y(P15[2]) );
  XNOR2X1 U263 ( .A(n67), .B(n36), .Y(P11[3]) );
  XOR2X1 U264 ( .A(P13[10]), .B(n24), .Y(P9[2]) );
  XOR2X1 U265 ( .A(n33), .B(n44), .Y(P7[2]) );
  XOR2X1 U266 ( .A(n45), .B(n46), .Y(P7[1]) );
  BUFX3 U267 ( .A(P3[4]), .Y(P4[8]) );
  XNOR2X1 U268 ( .A(n68), .B(P1[10]), .Y(n108) );
  CLKBUFXL U269 ( .A(P2[0]), .Y(P1[9]) );
  BUFX3 U270 ( .A(P2[11]), .Y(P1[7]) );
  XOR2X1 U271 ( .A(b_12), .B(P2[12]), .Y(n126) );
  XOR2X1 U272 ( .A(n3), .B(P1[10]), .Y(n127) );
  XNOR2X1 U273 ( .A(n88), .B(n89), .Y(n63) );
  XOR2X1 U274 ( .A(P6[11]), .B(n54), .Y(n44) );
  XNOR2X1 U275 ( .A(n128), .B(n129), .Y(n80) );
  XOR2X1 U276 ( .A(n19), .B(n78), .Y(n129) );
  BUFX3 U277 ( .A(b[8]), .Y(P1[12]) );
  XOR2X1 U278 ( .A(n130), .B(n131), .Y(P14[3]) );
  XOR2X1 U279 ( .A(n3), .B(n222), .Y(n130) );
  BUFX3 U280 ( .A(P5[10]), .Y(P4[6]) );
  XNOR2X1 U281 ( .A(n68), .B(P11[1]), .Y(P5[10]) );
  BUFX3 U282 ( .A(P6[0]), .Y(P5[9]) );
  BUFX3 U283 ( .A(P6[0]), .Y(P4[5]) );
  BUFX3 U284 ( .A(P6[12]), .Y(P4[4]) );
  XNOR2X1 U285 ( .A(n55), .B(n70), .Y(P6[12]) );
  BUFX3 U286 ( .A(P6[11]), .Y(P5[7]) );
  XOR2X1 U287 ( .A(P2[0]), .B(P12[2]), .Y(P6[11]) );
  BUFX3 U288 ( .A(P6[10]), .Y(P5[6]) );
  XNOR2X1 U289 ( .A(n61), .B(P12[1]), .Y(P6[10]) );
  BUFX3 U290 ( .A(P5[5]), .Y(P7[0]) );
  BUFX3 U291 ( .A(P5[5]), .Y(P6[9]) );
  BUFX3 U292 ( .A(P7[10]), .Y(P6[6]) );
  BUFX3 U293 ( .A(P7[7]), .Y(P8[11]) );
  XOR2X1 U294 ( .A(P3[10]), .B(n38), .Y(P7[7]) );
  BUFX3 U295 ( .A(P8[10]), .Y(P7[6]) );
  XNOR2X1 U296 ( .A(P1[10]), .B(n39), .Y(P8[10]) );
  BUFX3 U297 ( .A(P9[0]), .Y(P8[9]) );
  BUFX3 U298 ( .A(P9[0]), .Y(P7[5]) );
  BUFX3 U299 ( .A(P9[12]), .Y(P7[4]) );
  BUFX2 U300 ( .A(P9[11]), .Y(P8[7]) );
  XNOR2X1 U301 ( .A(n26), .B(n27), .Y(P9[11]) );
  BUFX3 U302 ( .A(P9[10]), .Y(P8[6]) );
  BUFX3 U303 ( .A(P9[9]), .Y(P10[0]) );
  BUFX3 U304 ( .A(P9[9]), .Y(P8[5]) );
  XNOR2XL U305 ( .A(n8), .B(P2[0]), .Y(n46) );
  XOR2X1 U306 ( .A(n91), .B(P2[10]), .Y(n97) );
  XNOR2X1 U307 ( .A(n67), .B(P2[0]), .Y(n86) );
  XNOR2XL U308 ( .A(n222), .B(b_12), .Y(n118) );
  XNOR2X1 U309 ( .A(n35), .B(n36), .Y(P8[2]) );
  XOR2X1 U310 ( .A(n120), .B(n123), .Y(P12[12]) );
  XNOR2X1 U311 ( .A(b[1]), .B(n34), .Y(P3[4]) );
  XNOR2XL U312 ( .A(n35), .B(n112), .Y(P3[1]) );
  XNOR2X1 U313 ( .A(b[1]), .B(n55), .Y(n114) );
  XNOR2XL U314 ( .A(n35), .B(n3), .Y(n84) );
  XNOR2X1 U315 ( .A(n35), .B(n68), .Y(n25) );
  XNOR2X1 U316 ( .A(n35), .B(P2[12]), .Y(n78) );
  XNOR2X1 U317 ( .A(P2[0]), .B(n35), .Y(n91) );
  XNOR2X1 U318 ( .A(n35), .B(b[3]), .Y(n53) );
  XNOR2X1 U319 ( .A(n3), .B(n56), .Y(n77) );
  XOR2X1 U320 ( .A(n53), .B(n44), .Y(P6[3]) );
  XNOR2X1 U321 ( .A(b[3]), .B(n34), .Y(P8[3]) );
  XNOR2X1 U322 ( .A(n67), .B(P11[2]), .Y(P4[7]) );
  XNOR2X1 U323 ( .A(n82), .B(P11[2]), .Y(P15[7]) );
  XOR2X1 U324 ( .A(n41), .B(n77), .Y(n122) );
  XOR2X1 U325 ( .A(n222), .B(n41), .Y(n120) );
  XOR2X1 U326 ( .A(b[3]), .B(P2[12]), .Y(n110) );
  XNOR2X1 U327 ( .A(n26), .B(b[3]), .Y(n111) );
  XNOR2X1 U328 ( .A(n56), .B(n17), .Y(P6[2]) );
  XNOR2X1 U329 ( .A(n56), .B(n76), .Y(P16[7]) );
  XNOR2X1 U330 ( .A(n56), .B(n110), .Y(n92) );
  XNOR2X1 U331 ( .A(n56), .B(n111), .Y(P3[2]) );
  XNOR2X1 U332 ( .A(n56), .B(n21), .Y(P12[2]) );
  XNOR2XL U333 ( .A(n55), .B(n1), .Y(n54) );
  XOR2X1 U334 ( .A(b_10), .B(n222), .Y(n59) );
  XOR2X1 U335 ( .A(b_10), .B(b[9]), .Y(P1[1]) );
  XNOR2XL U336 ( .A(n67), .B(n3), .Y(n24) );
  XNOR2X1 U337 ( .A(n3), .B(P1[12]), .Y(n57) );
  INVX8 U338 ( .A(b_11), .Y(n56) );
endmodule


module multiplier_column3_p16 ( b, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, 
        P11, P12, P13, P14, P15, P16 );
  input [12:0] b;
  output [12:0] P1;
  output [12:0] P2;
  output [12:0] P3;
  output [12:0] P4;
  output [12:0] P5;
  output [12:0] P6;
  output [12:0] P7;
  output [12:0] P8;
  output [12:0] P9;
  output [12:0] P10;
  output [12:0] P11;
  output [12:0] P12;
  output [12:0] P13;
  output [12:0] P14;
  output [12:0] P15;
  output [12:0] P16;
  wire   b_12, b_11, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n26,
         n27, n30, n31, n32, n33, n34, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n56, n57, n58,
         n60, n61, n62, n63, n64, n65, n66, n68, n69, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n84, n85, n86, n88, n89, n90, n91, n92,
         n94, n98, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n25, n28,
         n29, n35, n55, n59, n67, n70, n82, n83, n110, n174;
  assign b_12 = b[12];
  assign b_11 = b[11];

  XNOR2X1 U1 ( .A(n50), .B(P3[0]), .Y(n86) );
  INVX4 U2 ( .A(b[10]), .Y(n45) );
  XNOR2X1 U3 ( .A(n46), .B(n44), .Y(P6[0]) );
  XNOR2X2 U4 ( .A(n28), .B(P1[1]), .Y(P5[2]) );
  INVX1 U5 ( .A(b_11), .Y(n50) );
  XNOR2X2 U6 ( .A(P5[1]), .B(b[1]), .Y(n27) );
  XOR2X2 U7 ( .A(b[7]), .B(P1[11]), .Y(P2[1]) );
  OR2X2 U8 ( .A(n18), .B(n78), .Y(n10) );
  XOR2X1 U9 ( .A(n57), .B(n77), .Y(P13[9]) );
  OAI21XL U10 ( .A0(n40), .A1(n41), .B0(n8), .Y(n74) );
  NAND2X2 U11 ( .A(n9), .B(n10), .Y(n77) );
  XNOR2XL U12 ( .A(n45), .B(b[0]), .Y(n54) );
  INVX2 U13 ( .A(b[1]), .Y(n56) );
  XNOR2X2 U14 ( .A(n37), .B(n27), .Y(P8[7]) );
  NAND2X1 U15 ( .A(n6), .B(n7), .Y(n84) );
  NAND2X1 U16 ( .A(n4), .B(n5), .Y(n7) );
  XNOR2X1 U17 ( .A(n33), .B(n56), .Y(n30) );
  XOR2X1 U18 ( .A(P4[0]), .B(n90), .Y(n75) );
  XNOR2X2 U19 ( .A(P6[1]), .B(P2[11]), .Y(n18) );
  XOR2X1 U20 ( .A(P7[1]), .B(n59), .Y(P11[8]) );
  XNOR2X1 U21 ( .A(P2[3]), .B(n43), .Y(P5[1]) );
  CLKBUFX8 U22 ( .A(b[8]), .Y(P1[11]) );
  XNOR2X2 U23 ( .A(P3[3]), .B(n51), .Y(P6[1]) );
  BUFX3 U24 ( .A(P9[9]), .Y(P8[6]) );
  XNOR2X1 U25 ( .A(P4[3]), .B(n26), .Y(P7[1]) );
  XOR2X1 U26 ( .A(b_11), .B(n21), .Y(P16[2]) );
  BUFX3 U27 ( .A(P9[9]), .Y(P10[12]) );
  XNOR2XL U28 ( .A(b[3]), .B(n79), .Y(n62) );
  XOR2X2 U29 ( .A(b[6]), .B(P5[2]), .Y(n81) );
  XOR2X2 U30 ( .A(b[7]), .B(P3[0]), .Y(n39) );
  CLKBUFX3 U31 ( .A(P1[5]), .Y(P3[11]) );
  CLKBUFX3 U32 ( .A(P1[5]), .Y(P2[8]) );
  XOR2XL U33 ( .A(P2[0]), .B(n74), .Y(P11[2]) );
  XOR2X4 U34 ( .A(n81), .B(n89), .Y(P9[9]) );
  XNOR2X1 U35 ( .A(n51), .B(b[2]), .Y(n89) );
  XNOR2XL U36 ( .A(n51), .B(b[0]), .Y(n48) );
  INVX4 U37 ( .A(b[9]), .Y(n51) );
  XNOR2X2 U38 ( .A(n26), .B(b[5]), .Y(P3[2]) );
  XNOR2X1 U39 ( .A(b[10]), .B(n26), .Y(n15) );
  INVX4 U40 ( .A(b[6]), .Y(n26) );
  XNOR2XL U41 ( .A(n33), .B(b[5]), .Y(n91) );
  INVX2 U42 ( .A(b[3]), .Y(n33) );
  XNOR2X4 U43 ( .A(n45), .B(b_11), .Y(P1[1]) );
  XOR2X1 U44 ( .A(n72), .B(n75), .Y(P16[0]) );
  BUFX3 U45 ( .A(P16[0]), .Y(P13[4]) );
  INVX1 U46 ( .A(n86), .Y(n5) );
  INVX2 U47 ( .A(b[0]), .Y(n79) );
  INVX1 U48 ( .A(P3[0]), .Y(n44) );
  INVX4 U49 ( .A(b_12), .Y(n43) );
  XOR2X1 U50 ( .A(n19), .B(n20), .Y(P9[4]) );
  XNOR2X1 U51 ( .A(b[2]), .B(n52), .Y(P1[5]) );
  NAND2X1 U52 ( .A(n40), .B(n41), .Y(n8) );
  XNOR2X1 U53 ( .A(n34), .B(n43), .Y(P5[3]) );
  XOR2X1 U54 ( .A(n73), .B(n74), .Y(P15[11]) );
  XOR2X1 U55 ( .A(b[10]), .B(n53), .Y(P2[3]) );
  XNOR2X1 U56 ( .A(P1[11]), .B(b[0]), .Y(n28) );
  XOR2X1 U57 ( .A(b[1]), .B(P1[1]), .Y(P4[0]) );
  XNOR2X1 U58 ( .A(P6[0]), .B(n79), .Y(P13[1]) );
  BUFX3 U59 ( .A(P16[11]), .Y(P15[8]) );
  XOR2X1 U60 ( .A(n54), .B(n63), .Y(P16[12]) );
  XOR2X1 U61 ( .A(P2[0]), .B(n88), .Y(P13[10]) );
  BUFX3 U62 ( .A(b[7]), .Y(P2[0]) );
  CLKBUFX3 U63 ( .A(P13[11]), .Y(P11[5]) );
  XNOR2X1 U64 ( .A(n80), .B(n84), .Y(P13[11]) );
  XOR2XL U65 ( .A(n62), .B(n57), .Y(P15[2]) );
  XOR2XL U66 ( .A(b_12), .B(n57), .Y(n17) );
  BUFX2 U67 ( .A(P9[11]), .Y(P8[8]) );
  BUFX2 U68 ( .A(P9[11]), .Y(P7[5]) );
  XNOR2X2 U69 ( .A(n26), .B(n39), .Y(P3[3]) );
  XOR2X4 U70 ( .A(P9[9]), .B(n91), .Y(n88) );
  XNOR2XL U71 ( .A(n56), .B(n81), .Y(P12[3]) );
  BUFX3 U72 ( .A(b[5]), .Y(P2[11]) );
  XNOR2X1 U73 ( .A(P1[5]), .B(P2[11]), .Y(n40) );
  XNOR2X1 U74 ( .A(P1[11]), .B(P2[11]), .Y(n25) );
  XNOR2X1 U75 ( .A(b[2]), .B(P2[11]), .Y(n85) );
  XOR2X1 U76 ( .A(P16[2]), .B(P2[11]), .Y(P8[11]) );
  XOR2X1 U77 ( .A(b[5]), .B(P2[1]), .Y(n46) );
  XOR2X2 U78 ( .A(P2[1]), .B(n76), .Y(n65) );
  XNOR2X2 U79 ( .A(n79), .B(b[1]), .Y(n76) );
  NAND2XL U80 ( .A(P5[3]), .B(n86), .Y(n6) );
  INVX1 U81 ( .A(P5[3]), .Y(n4) );
  XNOR2X2 U82 ( .A(n33), .B(b_12), .Y(P2[9]) );
  BUFX1 U83 ( .A(P5[7]), .Y(P6[10]) );
  CLKBUFX2 U84 ( .A(P15[11]), .Y(P13[5]) );
  CLKBUFXL U85 ( .A(b[6]), .Y(P1[9]) );
  CLKBUFXL U86 ( .A(b[6]), .Y(P2[12]) );
  XNOR2XL U87 ( .A(n49), .B(b[1]), .Y(n78) );
  NAND2X1 U88 ( .A(n18), .B(n78), .Y(n9) );
  XOR2XL U89 ( .A(b[1]), .B(P3[1]), .Y(n12) );
  BUFX1 U90 ( .A(P12[12]), .Y(P10[6]) );
  XOR2X1 U91 ( .A(n72), .B(P10[3]), .Y(P13[6]) );
  BUFX1 U92 ( .A(P5[7]), .Y(P4[4]) );
  XNOR2X1 U93 ( .A(n26), .B(n75), .Y(P11[1]) );
  XNOR2X1 U94 ( .A(n44), .B(b[5]), .Y(P3[1]) );
  BUFX1 U95 ( .A(P13[6]), .Y(P15[12]) );
  XNOR2X1 U96 ( .A(n56), .B(n89), .Y(P15[1]) );
  CLKBUFXL U97 ( .A(P8[7]), .Y(P7[4]) );
  BUFX3 U98 ( .A(P6[11]), .Y(P5[8]) );
  BUFX3 U99 ( .A(P11[8]), .Y(P12[11]) );
  BUFX3 U100 ( .A(P13[11]), .Y(P12[8]) );
  XNOR2X1 U101 ( .A(n43), .B(P2[11]), .Y(n13) );
  XNOR2X1 U102 ( .A(n43), .B(b[1]), .Y(n94) );
  XOR2XL U103 ( .A(n26), .B(P3[0]), .Y(n14) );
  XOR2XL U104 ( .A(b[2]), .B(n53), .Y(n59) );
  XOR2X1 U105 ( .A(n82), .B(n57), .Y(n92) );
  XNOR2X1 U106 ( .A(b[0]), .B(P2[11]), .Y(n55) );
  BUFX8 U107 ( .A(b[4]), .Y(P3[0]) );
  CLKBUFXL U108 ( .A(P13[9]), .Y(P14[12]) );
  XOR2XL U109 ( .A(P2[2]), .B(P3[2]), .Y(P5[11]) );
  XNOR2XL U110 ( .A(P2[2]), .B(n52), .Y(P2[5]) );
  XNOR2X1 U111 ( .A(n39), .B(n40), .Y(P7[2]) );
  XNOR2XL U112 ( .A(n24), .B(n30), .Y(P8[3]) );
  XOR2X1 U113 ( .A(n21), .B(P16[3]), .Y(P12[12]) );
  BUFX2 U114 ( .A(P11[11]), .Y(P9[5]) );
  BUFX2 U115 ( .A(P11[11]), .Y(P10[8]) );
  CLKBUFXL U116 ( .A(P10[4]), .Y(P13[0]) );
  CLKBUFXL U117 ( .A(P10[4]), .Y(P11[7]) );
  CLKBUFXL U118 ( .A(P11[6]), .Y(P13[12]) );
  XNOR2XL U119 ( .A(n33), .B(b[2]), .Y(n72) );
  XNOR2X1 U120 ( .A(n26), .B(P2[3]), .Y(P3[6]) );
  XOR2X1 U121 ( .A(n20), .B(b[7]), .Y(n60) );
  XOR2X1 U122 ( .A(n11), .B(n61), .Y(P16[6]) );
  XOR2X1 U123 ( .A(P3[0]), .B(P2[9]), .Y(n11) );
  XNOR2X1 U124 ( .A(b[7]), .B(n51), .Y(n53) );
  XNOR2XL U125 ( .A(n17), .B(n18), .Y(P11[11]) );
  XOR2X1 U126 ( .A(n12), .B(n66), .Y(P14[1]) );
  XNOR2X1 U127 ( .A(n51), .B(n13), .Y(n36) );
  INVXL U128 ( .A(b[2]), .Y(n71) );
  XOR2X1 U129 ( .A(P1[2]), .B(n92), .Y(P9[11]) );
  XOR2X1 U130 ( .A(n88), .B(n94), .Y(P10[4]) );
  XOR2X1 U131 ( .A(n60), .B(n70), .Y(P10[3]) );
  XOR2XL U132 ( .A(n43), .B(P3[0]), .Y(n70) );
  XOR2X1 U133 ( .A(n84), .B(n85), .Y(P11[6]) );
  XNOR2X1 U134 ( .A(n24), .B(n14), .Y(P9[1]) );
  XNOR2X1 U135 ( .A(n26), .B(b[1]), .Y(n58) );
  XNOR2X1 U136 ( .A(b[2]), .B(n19), .Y(P12[2]) );
  XNOR2X1 U137 ( .A(n45), .B(n46), .Y(P6[2]) );
  XOR2X1 U138 ( .A(n62), .B(n77), .Y(P12[5]) );
  XOR2XL U139 ( .A(P1[11]), .B(P3[0]), .Y(n82) );
  XOR2X1 U140 ( .A(n27), .B(n25), .Y(P8[5]) );
  INVX1 U141 ( .A(P1[2]), .Y(n52) );
  XNOR2XL U142 ( .A(b[3]), .B(n50), .Y(n37) );
  XNOR2XL U143 ( .A(b[3]), .B(n26), .Y(n80) );
  XNOR2XL U144 ( .A(n68), .B(b_11), .Y(n32) );
  XNOR2X1 U145 ( .A(b_11), .B(n43), .Y(P1[2]) );
  XNOR2X1 U146 ( .A(P4[1]), .B(n29), .Y(P16[4]) );
  XOR2X1 U147 ( .A(n26), .B(b[9]), .Y(n29) );
  XOR2XL U148 ( .A(b[9]), .B(n92), .Y(n68) );
  XOR2X1 U149 ( .A(n35), .B(n65), .Y(n34) );
  XOR2X1 U150 ( .A(b[10]), .B(b[9]), .Y(n35) );
  XOR2X1 U151 ( .A(n32), .B(n55), .Y(P14[3]) );
  BUFX3 U152 ( .A(P5[11]), .Y(P3[5]) );
  CLKBUFXL U153 ( .A(P16[0]), .Y(P14[7]) );
  CLKBUFXL U154 ( .A(P16[0]), .Y(P15[10]) );
  BUFX3 U155 ( .A(P9[0]), .Y(P8[10]) );
  BUFX3 U156 ( .A(P9[0]), .Y(P6[4]) );
  INVX1 U157 ( .A(P13[7]), .Y(n110) );
  INVXL U158 ( .A(P6[0]), .Y(n174) );
  BUFX3 U159 ( .A(P2[5]), .Y(P4[11]) );
  BUFX3 U160 ( .A(P2[5]), .Y(P3[8]) );
  CLKBUFXL U161 ( .A(P13[9]), .Y(P12[6]) );
  BUFX3 U162 ( .A(P12[12]), .Y(P11[9]) );
  BUFX3 U163 ( .A(P13[6]), .Y(P14[9]) );
  BUFX3 U164 ( .A(P5[11]), .Y(P4[8]) );
  XNOR2X1 U165 ( .A(n44), .B(P16[1]), .Y(P9[0]) );
  XNOR2X1 U166 ( .A(n44), .B(n36), .Y(P16[7]) );
  XOR2X1 U167 ( .A(P9[11]), .B(n91), .Y(P16[3]) );
  XNOR2X1 U168 ( .A(n49), .B(P15[2]), .Y(P7[11]) );
  BUFX3 U169 ( .A(P7[11]), .Y(P6[8]) );
  XNOR2X1 U170 ( .A(n44), .B(n64), .Y(n38) );
  XNOR2X1 U171 ( .A(n30), .B(n86), .Y(n47) );
  XNOR2X1 U172 ( .A(n21), .B(n22), .Y(P9[3]) );
  XNOR2X1 U173 ( .A(n22), .B(n91), .Y(P10[2]) );
  XOR2X1 U174 ( .A(n53), .B(n38), .Y(P10[1]) );
  INVX1 U175 ( .A(n110), .Y(P12[4]) );
  INVXL U176 ( .A(n110), .Y(P14[10]) );
  XOR2X1 U177 ( .A(P16[5]), .B(n78), .Y(P12[1]) );
  BUFX3 U178 ( .A(P16[7]), .Y(P15[4]) );
  BUFX3 U179 ( .A(P16[8]), .Y(P15[5]) );
  BUFX3 U180 ( .A(P9[12]), .Y(P7[6]) );
  BUFX3 U181 ( .A(P9[0]), .Y(P7[7]) );
  BUFX3 U182 ( .A(P7[11]), .Y(P5[5]) );
  BUFX3 U183 ( .A(P6[12]), .Y(P5[9]) );
  BUFX3 U184 ( .A(P3[7]), .Y(P4[10]) );
  BUFX3 U185 ( .A(P5[7]), .Y(P7[0]) );
  BUFX3 U186 ( .A(P6[11]), .Y(P4[5]) );
  BUFX3 U187 ( .A(P5[4]), .Y(P8[0]) );
  BUFX3 U188 ( .A(P3[7]), .Y(P5[0]) );
  BUFX3 U189 ( .A(P3[7]), .Y(P2[4]) );
  BUFX3 U190 ( .A(P15[7]), .Y(P16[10]) );
  CLKBUFXL U191 ( .A(P4[0]), .Y(P3[10]) );
  CLKBUFXL U192 ( .A(P4[0]), .Y(P2[7]) );
  CLKBUFXL U193 ( .A(P4[0]), .Y(P1[4]) );
  BUFX3 U194 ( .A(P9[4]), .Y(P12[0]) );
  BUFX3 U195 ( .A(P9[4]), .Y(P11[10]) );
  BUFX3 U196 ( .A(P9[4]), .Y(P10[7]) );
  CLKBUFXL U197 ( .A(P10[4]), .Y(P12[10]) );
  BUFX3 U198 ( .A(P15[6]), .Y(P16[9]) );
  BUFX3 U199 ( .A(P16[12]), .Y(P14[6]) );
  BUFX3 U200 ( .A(P16[12]), .Y(P15[9]) );
  BUFX3 U201 ( .A(P8[11]), .Y(P7[8]) );
  BUFX3 U202 ( .A(P8[11]), .Y(P6[5]) );
  BUFX3 U203 ( .A(P5[4]), .Y(P7[10]) );
  BUFX3 U204 ( .A(P6[6]), .Y(P8[12]) );
  BUFX3 U205 ( .A(P6[6]), .Y(P7[9]) );
  BUFX3 U206 ( .A(P12[5]), .Y(P14[11]) );
  BUFX3 U207 ( .A(P12[5]), .Y(P13[8]) );
  BUFX3 U208 ( .A(P11[8]), .Y(P10[5]) );
  BUFX3 U209 ( .A(P9[6]), .Y(P11[12]) );
  BUFX3 U210 ( .A(P9[6]), .Y(P10[9]) );
  BUFX3 U211 ( .A(P3[6]), .Y(P4[9]) );
  BUFX3 U212 ( .A(P3[9]), .Y(P2[6]) );
  BUFX3 U213 ( .A(P6[12]), .Y(P4[6]) );
  BUFX3 U214 ( .A(P8[5]), .Y(P9[8]) );
  BUFX3 U215 ( .A(P8[5]), .Y(P10[11]) );
  BUFX3 U216 ( .A(P11[6]), .Y(P12[9]) );
  BUFX3 U217 ( .A(P15[11]), .Y(P14[8]) );
  BUFX3 U218 ( .A(P16[11]), .Y(P14[5]) );
  BUFX3 U219 ( .A(P9[12]), .Y(P8[9]) );
  BUFX3 U220 ( .A(P7[12]), .Y(P6[9]) );
  BUFX3 U221 ( .A(P7[12]), .Y(P5[6]) );
  BUFX3 U222 ( .A(P8[7]), .Y(P9[10]) );
  CLKBUFXL U223 ( .A(P8[7]), .Y(P10[0]) );
  BUFX3 U224 ( .A(P13[10]), .Y(P11[4]) );
  BUFX3 U225 ( .A(P13[10]), .Y(P12[7]) );
  BUFX3 U226 ( .A(P13[10]), .Y(P14[0]) );
  BUFX3 U227 ( .A(P5[4]), .Y(P6[7]) );
  XNOR2X1 U228 ( .A(n45), .B(P14[1]), .Y(P5[7]) );
  XOR2X1 U229 ( .A(P2[0]), .B(P15[1]), .Y(P5[4]) );
  XNOR2X1 U230 ( .A(n45), .B(b[2]), .Y(n57) );
  INVX1 U231 ( .A(n174), .Y(P5[10]) );
  XNOR2X1 U232 ( .A(b[7]), .B(n79), .Y(n21) );
  XOR2X1 U233 ( .A(n41), .B(n42), .Y(P6[6]) );
  XNOR2XL U234 ( .A(n43), .B(P1[11]), .Y(n42) );
  XNOR2X1 U235 ( .A(n50), .B(P14[2]), .Y(P6[11]) );
  XNOR2X1 U236 ( .A(n51), .B(P1[3]), .Y(P3[9]) );
  XNOR2X1 U237 ( .A(n15), .B(n16), .Y(P9[6]) );
  XOR2X1 U238 ( .A(P3[3]), .B(P2[9]), .Y(P6[12]) );
  XOR2X1 U239 ( .A(n64), .B(n48), .Y(P16[11]) );
  XOR2X1 U240 ( .A(n37), .B(n36), .Y(P9[12]) );
  XOR2X1 U241 ( .A(P3[2]), .B(n54), .Y(P16[8]) );
  XNOR2X1 U242 ( .A(n43), .B(n15), .Y(P16[1]) );
  XOR2X1 U243 ( .A(n47), .B(n48), .Y(P7[12]) );
  XNOR2X1 U244 ( .A(P4[2]), .B(n67), .Y(P16[5]) );
  XOR2X1 U245 ( .A(P2[0]), .B(n45), .Y(n67) );
  XNOR2X1 U246 ( .A(P1[11]), .B(n51), .Y(P2[2]) );
  XOR2X1 U247 ( .A(P16[2]), .B(n58), .Y(P15[6]) );
  XNOR2X1 U248 ( .A(n43), .B(n54), .Y(P1[3]) );
  XNOR2X1 U249 ( .A(n46), .B(n37), .Y(n16) );
  XNOR2XL U250 ( .A(n69), .B(P2[11]), .Y(P14[2]) );
  XOR2X1 U251 ( .A(n73), .B(P15[1]), .Y(n63) );
  XNOR2X1 U252 ( .A(b[1]), .B(P3[2]), .Y(n20) );
  XNOR2X1 U253 ( .A(n30), .B(n98), .Y(n64) );
  XNOR2XL U254 ( .A(n71), .B(P1[11]), .Y(n98) );
  XNOR2X1 U255 ( .A(n56), .B(n17), .Y(P4[1]) );
  XOR2X1 U256 ( .A(n31), .B(n47), .Y(P4[3]) );
  XOR2X1 U257 ( .A(P8[11]), .B(n31), .Y(n24) );
  BUFX3 U258 ( .A(P15[7]), .Y(P14[4]) );
  XNOR2X1 U259 ( .A(n50), .B(n63), .Y(P11[3]) );
  XNOR2X1 U260 ( .A(b[1]), .B(n32), .Y(P8[2]) );
  XNOR2X1 U261 ( .A(b[2]), .B(n23), .Y(P15[3]) );
  XNOR2XL U262 ( .A(n33), .B(n34), .Y(P8[1]) );
  INVX1 U263 ( .A(n174), .Y(P4[7]) );
  INVX1 U264 ( .A(n174), .Y(P3[4]) );
  INVXL U265 ( .A(n110), .Y(P15[0]) );
  XOR2X1 U266 ( .A(n15), .B(n38), .Y(P7[3]) );
  XNOR2X1 U267 ( .A(b[2]), .B(n80), .Y(n69) );
  INVX1 U268 ( .A(n68), .Y(n22) );
  BUFX3 U269 ( .A(P2[9]), .Y(P3[12]) );
  BUFX3 U270 ( .A(P3[9]), .Y(P4[12]) );
  BUFX3 U271 ( .A(P3[6]), .Y(P5[12]) );
  INVXL U272 ( .A(P1[11]), .Y(n49) );
  BUFX3 U273 ( .A(P10[10]), .Y(P11[0]) );
  BUFX3 U274 ( .A(P10[10]), .Y(P9[7]) );
  BUFX3 U275 ( .A(P10[10]), .Y(P8[4]) );
  CLKBUFXL U276 ( .A(P2[0]), .Y(P1[10]) );
  CLKBUFXL U277 ( .A(P3[0]), .Y(P2[10]) );
  CLKBUFXL U278 ( .A(P3[0]), .Y(P1[7]) );
  BUFX3 U279 ( .A(P2[9]), .Y(P1[6]) );
  CLKBUFXL U280 ( .A(P2[11]), .Y(P1[8]) );
  XOR2X1 U281 ( .A(P2[5]), .B(n83), .Y(P10[10]) );
  XOR2X1 U282 ( .A(P3[3]), .B(b[0]), .Y(n83) );
  XNOR2X1 U283 ( .A(b[10]), .B(n43), .Y(n31) );
  XNOR2X1 U284 ( .A(P16[6]), .B(b[9]), .Y(n19) );
  XNOR2XL U285 ( .A(n71), .B(b_12), .Y(n66) );
  XNOR2X1 U286 ( .A(b[3]), .B(n44), .Y(n73) );
  XNOR2X1 U287 ( .A(b_12), .B(n23), .Y(P9[2]) );
  XNOR2X1 U288 ( .A(b_12), .B(n16), .Y(P13[3]) );
  CLKBUFXL U289 ( .A(b[9]), .Y(P1[12]) );
  CLKBUFXL U290 ( .A(b[10]), .Y(P1[0]) );
  XOR2X1 U291 ( .A(n76), .B(P5[11]), .Y(P13[2]) );
  XOR2X1 U292 ( .A(n65), .B(n66), .Y(P15[7]) );
  XNOR2X1 U293 ( .A(n69), .B(P13[1]), .Y(P13[7]) );
  XOR2X1 U294 ( .A(P2[1]), .B(P1[1]), .Y(P3[7]) );
  XNOR2X1 U295 ( .A(n79), .B(n58), .Y(n41) );
  XNOR2X1 U296 ( .A(n79), .B(P3[1]), .Y(n90) );
  XOR2X1 U297 ( .A(n60), .B(n61), .Y(n23) );
  XNOR2X1 U298 ( .A(n49), .B(b_11), .Y(n61) );
  XNOR2X1 U299 ( .A(b_11), .B(n18), .Y(P6[3]) );
  XOR2X1 U300 ( .A(b_11), .B(n72), .Y(P4[2]) );
endmodule


module multiplier_column2_p16 ( b, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, 
        P11, P12, P13, P14, P15, P16 );
  input [12:0] b;
  output [12:0] P1;
  output [12:0] P2;
  output [12:0] P3;
  output [12:0] P4;
  output [12:0] P5;
  output [12:0] P6;
  output [12:0] P7;
  output [12:0] P8;
  output [12:0] P9;
  output [12:0] P10;
  output [12:0] P11;
  output [12:0] P12;
  output [12:0] P13;
  output [12:0] P14;
  output [12:0] P15;
  output [12:0] P16;
  wire   b_12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n86,
         n87, n88, n89, n90, n91, n1, n3, n4, n5, n6, n205;
  assign b_12 = b[12];

  XNOR2X4 U19 ( .A(b[1]), .B(n34), .Y(P10[12]) );
  XNOR2X4 U42 ( .A(n1), .B(n40), .Y(n34) );
  XNOR2X4 U78 ( .A(n53), .B(b[6]), .Y(P4[2]) );
  XOR2X4 U85 ( .A(n75), .B(n76), .Y(P13[7]) );
  XOR2X4 U103 ( .A(n75), .B(n80), .Y(P15[0]) );
  XNOR2X4 U105 ( .A(P8[2]), .B(b[1]), .Y(n75) );
  BUFX4 U1 ( .A(b[7]), .Y(P3[0]) );
  XNOR2X1 U2 ( .A(n56), .B(n19), .Y(n67) );
  XNOR2X2 U3 ( .A(n39), .B(n40), .Y(n56) );
  XOR2X2 U4 ( .A(b[0]), .B(b[11]), .Y(n66) );
  XNOR2X4 U5 ( .A(n71), .B(n38), .Y(n39) );
  XNOR2X4 U6 ( .A(b_12), .B(P4[2]), .Y(n71) );
  INVX4 U7 ( .A(P3[0]), .Y(n53) );
  XNOR2X1 U8 ( .A(n41), .B(n66), .Y(n33) );
  XNOR2X1 U9 ( .A(n37), .B(P4[12]), .Y(n1) );
  CLKINVX3 U10 ( .A(b[10]), .Y(n19) );
  XNOR2X2 U11 ( .A(b[9]), .B(n41), .Y(P3[2]) );
  XNOR2XL U12 ( .A(b[2]), .B(n41), .Y(n57) );
  INVX2 U13 ( .A(b[8]), .Y(n41) );
  XOR2X1 U14 ( .A(n46), .B(n5), .Y(n43) );
  XNOR2X2 U15 ( .A(n54), .B(n67), .Y(P16[10]) );
  XNOR2X1 U16 ( .A(b[2]), .B(n19), .Y(n82) );
  XOR2XL U17 ( .A(b[2]), .B(b[9]), .Y(n54) );
  XOR2X1 U18 ( .A(P6[3]), .B(P2[10]), .Y(P11[2]) );
  XOR2X1 U20 ( .A(b_12), .B(n82), .Y(n37) );
  BUFX3 U21 ( .A(b[4]), .Y(P4[12]) );
  XNOR2X2 U22 ( .A(P3[3]), .B(n31), .Y(P8[2]) );
  CLKINVX3 U23 ( .A(b_12), .Y(n31) );
  XOR2X1 U24 ( .A(n79), .B(n81), .Y(P14[10]) );
  XOR2X1 U25 ( .A(n63), .B(n64), .Y(P16[8]) );
  BUFX3 U26 ( .A(P16[10]), .Y(P13[4]) );
  XNOR2XL U27 ( .A(n73), .B(P3[0]), .Y(n77) );
  XNOR2XL U28 ( .A(n31), .B(P3[0]), .Y(n91) );
  XNOR2XL U29 ( .A(n42), .B(P3[0]), .Y(n13) );
  XNOR2XL U30 ( .A(n78), .B(P3[0]), .Y(n63) );
  XNOR2X1 U31 ( .A(P3[0]), .B(n62), .Y(P13[1]) );
  XOR2X2 U32 ( .A(P1[1]), .B(n30), .Y(n86) );
  XNOR2X2 U33 ( .A(n19), .B(n205), .Y(n30) );
  BUFX2 U34 ( .A(P16[8]), .Y(P15[6]) );
  BUFX3 U35 ( .A(P16[8]), .Y(P14[4]) );
  BUFX3 U36 ( .A(b[6]), .Y(P2[10]) );
  XNOR2X1 U37 ( .A(n23), .B(n14), .Y(n62) );
  XNOR2X1 U38 ( .A(n40), .B(P4[12]), .Y(P5[2]) );
  XNOR2X1 U39 ( .A(n33), .B(n77), .Y(n24) );
  XNOR2XL U40 ( .A(P2[10]), .B(n24), .Y(P8[3]) );
  CLKBUFX2 U41 ( .A(P14[5]), .Y(P15[7]) );
  XOR2X1 U43 ( .A(n22), .B(P11[2]), .Y(P16[7]) );
  CLKBUFX2 U44 ( .A(P13[7]), .Y(P16[0]) );
  XNOR2X2 U45 ( .A(n73), .B(b[10]), .Y(P2[1]) );
  XOR2X1 U46 ( .A(P2[9]), .B(b[10]), .Y(n3) );
  BUFX3 U47 ( .A(P16[7]), .Y(P15[5]) );
  BUFX2 U48 ( .A(P4[7]), .Y(P5[9]) );
  BUFX2 U49 ( .A(P4[7]), .Y(P3[5]) );
  BUFX1 U50 ( .A(P4[7]), .Y(P6[11]) );
  XNOR2XL U51 ( .A(n41), .B(P3[0]), .Y(P3[1]) );
  XOR2X1 U52 ( .A(n43), .B(n45), .Y(P16[4]) );
  XNOR2X2 U53 ( .A(b[11]), .B(n31), .Y(P1[1]) );
  XNOR2X1 U54 ( .A(P4[12]), .B(b[1]), .Y(n4) );
  XNOR2X1 U55 ( .A(b[9]), .B(b[0]), .Y(n32) );
  XOR2XL U56 ( .A(n21), .B(b[10]), .Y(n5) );
  CLKBUFXL U57 ( .A(P13[5]), .Y(P14[7]) );
  CLKBUFXL U58 ( .A(P13[5]), .Y(P15[9]) );
  XOR2XL U59 ( .A(n29), .B(n30), .Y(P7[4]) );
  XOR2XL U60 ( .A(P6[2]), .B(P4[1]), .Y(P9[11]) );
  XNOR2X1 U61 ( .A(n61), .B(n62), .Y(P14[5]) );
  BUFX3 U62 ( .A(P16[10]), .Y(P15[8]) );
  CLKINVX3 U63 ( .A(P2[9]), .Y(n40) );
  XNOR2XL U64 ( .A(n35), .B(n40), .Y(n14) );
  XNOR2XL U65 ( .A(n31), .B(n205), .Y(P1[5]) );
  INVXL U66 ( .A(n205), .Y(n28) );
  XNOR2XL U67 ( .A(n28), .B(P4[12]), .Y(n27) );
  XNOR2XL U68 ( .A(n73), .B(P1[1]), .Y(P2[3]) );
  XNOR2X1 U69 ( .A(n205), .B(n34), .Y(P16[3]) );
  XOR2X1 U70 ( .A(P3[0]), .B(P2[1]), .Y(P3[3]) );
  XNOR2XL U71 ( .A(n21), .B(n205), .Y(n50) );
  XNOR2XL U72 ( .A(n73), .B(n205), .Y(n69) );
  XNOR2XL U73 ( .A(n79), .B(n21), .Y(P7[3]) );
  XNOR2X1 U74 ( .A(n21), .B(n22), .Y(P11[11]) );
  XNOR2X1 U75 ( .A(P2[10]), .B(n46), .Y(P12[4]) );
  XOR2XL U76 ( .A(P3[2]), .B(P4[1]), .Y(P8[12]) );
  XNOR2X1 U77 ( .A(n55), .B(n31), .Y(n23) );
  XNOR2X1 U79 ( .A(n21), .B(n37), .Y(P6[1]) );
  CLKBUFXL U80 ( .A(P4[12]), .Y(P3[10]) );
  CLKBUFXL U81 ( .A(P2[9]), .Y(P3[11]) );
  CLKBUFXL U82 ( .A(P4[12]), .Y(P1[6]) );
  XNOR2XL U83 ( .A(n21), .B(n63), .Y(P12[3]) );
  XNOR2X1 U84 ( .A(n55), .B(P11[1]), .Y(P15[4]) );
  BUFX3 U86 ( .A(P10[12]), .Y(P9[10]) );
  CLKBUFXL U87 ( .A(P2[9]), .Y(P4[0]) );
  CLKBUFXL U88 ( .A(P4[12]), .Y(P2[8]) );
  CLKBUFXL U89 ( .A(P2[9]), .Y(P1[7]) );
  CLKINVX3 U90 ( .A(b[1]), .Y(n21) );
  XOR2XL U91 ( .A(b[2]), .B(P1[1]), .Y(P1[4]) );
  XNOR2XL U92 ( .A(n35), .B(b[1]), .Y(P1[3]) );
  INVX1 U93 ( .A(b[9]), .Y(n73) );
  XOR2X1 U94 ( .A(n3), .B(n61), .Y(n58) );
  XNOR2XL U95 ( .A(b[2]), .B(P2[9]), .Y(n44) );
  XNOR2XL U96 ( .A(n42), .B(b_12), .Y(P1[2]) );
  XNOR2XL U97 ( .A(b[0]), .B(b[1]), .Y(n83) );
  XNOR2XL U98 ( .A(b[0]), .B(n23), .Y(P12[12]) );
  XOR2X1 U99 ( .A(n1), .B(n89), .Y(P13[10]) );
  XOR2X1 U100 ( .A(b[8]), .B(n6), .Y(n55) );
  XNOR2X1 U101 ( .A(n4), .B(n86), .Y(P6[3]) );
  XNOR2XL U102 ( .A(b[8]), .B(P2[9]), .Y(n76) );
  XOR2X1 U104 ( .A(n87), .B(n86), .Y(n78) );
  XNOR2XL U106 ( .A(b[0]), .B(P2[9]), .Y(n87) );
  XNOR2XL U107 ( .A(b[11]), .B(n205), .Y(n80) );
  CLKBUFXL U108 ( .A(b[11]), .Y(P1[0]) );
  BUFX3 U109 ( .A(P13[0]), .Y(P12[11]) );
  BUFX3 U110 ( .A(P13[0]), .Y(P10[7]) );
  BUFX3 U111 ( .A(P13[0]), .Y(P9[5]) );
  BUFX3 U112 ( .A(P9[11]), .Y(P6[5]) );
  BUFX3 U113 ( .A(P7[4]), .Y(P8[6]) );
  BUFX3 U114 ( .A(P13[5]), .Y(P16[11]) );
  BUFX3 U115 ( .A(P6[7]), .Y(P8[11]) );
  BUFX3 U116 ( .A(P6[7]), .Y(P7[9]) );
  BUFX3 U117 ( .A(P7[11]), .Y(P6[9]) );
  BUFX3 U118 ( .A(P6[7]), .Y(P5[5]) );
  BUFX3 U119 ( .A(P7[11]), .Y(P5[7]) );
  BUFX3 U120 ( .A(P7[4]), .Y(P11[12]) );
  BUFX3 U121 ( .A(P7[4]), .Y(P10[10]) );
  BUFX3 U122 ( .A(P7[4]), .Y(P9[8]) );
  BUFX3 U123 ( .A(P9[11]), .Y(P10[0]) );
  BUFX3 U124 ( .A(P9[11]), .Y(P8[9]) );
  BUFX3 U125 ( .A(P9[11]), .Y(P7[7]) );
  BUFX3 U126 ( .A(P14[5]), .Y(P16[9]) );
  XNOR2X1 U127 ( .A(n13), .B(n14), .Y(P13[0]) );
  XNOR2X1 U128 ( .A(n17), .B(P3[3]), .Y(P7[11]) );
  XNOR2X1 U129 ( .A(n38), .B(P4[3]), .Y(P6[7]) );
  XOR2X1 U130 ( .A(n70), .B(P3[4]), .Y(P13[5]) );
  XNOR2X1 U131 ( .A(n40), .B(P3[1]), .Y(P4[3]) );
  XNOR2X1 U132 ( .A(n53), .B(n65), .Y(n60) );
  XNOR2X1 U133 ( .A(n38), .B(n77), .Y(n20) );
  XNOR2X1 U134 ( .A(n14), .B(n20), .Y(n18) );
  XOR2X1 U135 ( .A(n24), .B(n15), .Y(n46) );
  XOR2X1 U136 ( .A(n49), .B(n50), .Y(P16[2]) );
  BUFX3 U137 ( .A(P6[7]), .Y(P9[0]) );
  BUFX3 U138 ( .A(P8[12]), .Y(P6[8]) );
  BUFX3 U139 ( .A(P3[4]), .Y(P6[10]) );
  BUFX3 U140 ( .A(P7[11]), .Y(P4[5]) );
  BUFX3 U141 ( .A(P11[11]), .Y(P9[7]) );
  XNOR2X1 U142 ( .A(n17), .B(n25), .Y(P8[1]) );
  BUFX3 U143 ( .A(P11[11]), .Y(P8[5]) );
  BUFX3 U144 ( .A(P10[5]), .Y(P12[9]) );
  BUFX3 U145 ( .A(P13[0]), .Y(P11[9]) );
  BUFX3 U146 ( .A(P11[11]), .Y(P10[9]) );
  XOR2X1 U147 ( .A(n13), .B(n72), .Y(P12[1]) );
  XNOR2X1 U148 ( .A(n17), .B(n18), .Y(P9[3]) );
  BUFX3 U149 ( .A(P9[9]), .Y(P7[5]) );
  BUFX3 U150 ( .A(P8[12]), .Y(P4[4]) );
  BUFX3 U151 ( .A(P10[5]), .Y(P13[11]) );
  XNOR2XL U152 ( .A(n14), .B(n72), .Y(P13[3]) );
  XNOR2X1 U153 ( .A(n38), .B(P1[5]), .Y(P5[1]) );
  XNOR2X1 U154 ( .A(n17), .B(n20), .Y(P9[1]) );
  XNOR2X1 U155 ( .A(n17), .B(n60), .Y(P14[3]) );
  BUFX3 U156 ( .A(P12[4]), .Y(P16[12]) );
  BUFX3 U157 ( .A(P3[4]), .Y(P5[8]) );
  BUFX3 U158 ( .A(P3[4]), .Y(P4[6]) );
  BUFX3 U159 ( .A(P12[4]), .Y(P14[8]) );
  BUFX3 U160 ( .A(P12[4]), .Y(P15[10]) );
  BUFX3 U161 ( .A(P12[4]), .Y(P13[6]) );
  BUFX3 U162 ( .A(P11[11]), .Y(P12[0]) );
  BUFX3 U163 ( .A(P5[4]), .Y(P8[10]) );
  BUFX3 U164 ( .A(P5[4]), .Y(P7[8]) );
  BUFX3 U165 ( .A(P5[4]), .Y(P6[6]) );
  BUFX3 U166 ( .A(P6[0]), .Y(P5[11]) );
  BUFX3 U167 ( .A(P6[0]), .Y(P4[9]) );
  BUFX3 U168 ( .A(P6[0]), .Y(P2[5]) );
  BUFX3 U169 ( .A(P6[0]), .Y(P3[7]) );
  BUFX3 U170 ( .A(P8[12]), .Y(P7[10]) );
  BUFX3 U171 ( .A(P8[12]), .Y(P5[6]) );
  BUFX3 U172 ( .A(P10[5]), .Y(P11[7]) );
  BUFX3 U173 ( .A(P5[10]), .Y(P4[8]) );
  BUFX3 U174 ( .A(P5[10]), .Y(P2[4]) );
  BUFX3 U175 ( .A(P10[5]), .Y(P14[0]) );
  BUFX3 U176 ( .A(P9[9]), .Y(P11[0]) );
  BUFX3 U177 ( .A(P9[9]), .Y(P10[11]) );
  BUFX3 U178 ( .A(P9[9]), .Y(P8[7]) );
  BUFX3 U179 ( .A(P14[10]), .Y(P12[6]) );
  BUFX3 U180 ( .A(P14[10]), .Y(P11[4]) );
  BUFX3 U181 ( .A(P14[10]), .Y(P15[12]) );
  BUFX3 U182 ( .A(P14[10]), .Y(P13[8]) );
  BUFX3 U183 ( .A(P16[10]), .Y(P14[6]) );
  BUFX3 U184 ( .A(P15[4]), .Y(P16[6]) );
  BUFX3 U185 ( .A(P1[5]), .Y(P5[0]) );
  BUFX3 U186 ( .A(P1[5]), .Y(P4[11]) );
  BUFX3 U187 ( .A(P1[5]), .Y(P2[7]) );
  INVX1 U188 ( .A(n53), .Y(P1[9]) );
  XOR2X1 U189 ( .A(P2[2]), .B(P3[1]), .Y(P3[4]) );
  XNOR2X1 U190 ( .A(n41), .B(P2[3]), .Y(P4[7]) );
  XNOR2X1 U191 ( .A(n19), .B(P1[3]), .Y(P6[0]) );
  XNOR2X1 U192 ( .A(n205), .B(n39), .Y(P5[4]) );
  XOR2X1 U193 ( .A(P2[1]), .B(P1[2]), .Y(P5[10]) );
  XOR2X1 U194 ( .A(P2[3]), .B(n88), .Y(P10[5]) );
  XNOR2XL U195 ( .A(n28), .B(P2[9]), .Y(n88) );
  XOR2X1 U196 ( .A(n26), .B(n27), .Y(P9[9]) );
  XNOR2XL U197 ( .A(n42), .B(P2[10]), .Y(n81) );
  XNOR2X1 U198 ( .A(n40), .B(P1[8]), .Y(P4[1]) );
  XNOR2X1 U199 ( .A(n41), .B(n59), .Y(n64) );
  INVX1 U200 ( .A(P4[12]), .Y(n38) );
  XNOR2X1 U201 ( .A(n19), .B(n65), .Y(n72) );
  XOR2X1 U202 ( .A(P3[2]), .B(n50), .Y(n65) );
  XNOR2X1 U203 ( .A(n31), .B(P4[12]), .Y(n15) );
  XNOR2X1 U204 ( .A(n53), .B(n54), .Y(n22) );
  XNOR2X1 U205 ( .A(n71), .B(n29), .Y(n49) );
  XNOR2X1 U206 ( .A(n35), .B(P3[2]), .Y(n25) );
  XNOR2X1 U207 ( .A(n44), .B(n91), .Y(n84) );
  XNOR2X1 U208 ( .A(n42), .B(n57), .Y(n29) );
  XNOR2X1 U209 ( .A(n78), .B(n54), .Y(P11[1]) );
  XNOR2X1 U210 ( .A(n70), .B(n31), .Y(P5[3]) );
  XOR2X1 U211 ( .A(P4[12]), .B(n69), .Y(n61) );
  INVXL U212 ( .A(P2[10]), .Y(n17) );
  XNOR2X1 U213 ( .A(n43), .B(n44), .Y(P16[5]) );
  XOR2X1 U214 ( .A(n51), .B(n52), .Y(P16[1]) );
  XNOR2XL U215 ( .A(n28), .B(P2[10]), .Y(n45) );
  XNOR2X1 U216 ( .A(n35), .B(n36), .Y(P6[2]) );
  XOR2X1 U217 ( .A(n25), .B(n82), .Y(n79) );
  XOR2X1 U218 ( .A(n205), .B(P4[1]), .Y(n70) );
  BUFX3 U219 ( .A(P5[4]), .Y(P9[12]) );
  BUFX3 U220 ( .A(P7[11]), .Y(P8[0]) );
  BUFX3 U221 ( .A(P4[7]), .Y(P7[0]) );
  BUFX3 U222 ( .A(P3[4]), .Y(P7[12]) );
  BUFX3 U223 ( .A(P5[10]), .Y(P6[12]) );
  BUFX3 U224 ( .A(P1[4]), .Y(P5[12]) );
  BUFX3 U225 ( .A(P1[4]), .Y(P4[10]) );
  XNOR2X1 U226 ( .A(n41), .B(P5[3]), .Y(P10[2]) );
  BUFX3 U227 ( .A(P9[4]), .Y(P11[8]) );
  XNOR2XL U228 ( .A(n31), .B(n26), .Y(P7[2]) );
  XOR2X1 U229 ( .A(n57), .B(n58), .Y(P15[2]) );
  BUFX3 U230 ( .A(P9[4]), .Y(P12[10]) );
  BUFX3 U231 ( .A(P9[4]), .Y(P13[12]) );
  BUFX3 U232 ( .A(P9[4]), .Y(P10[6]) );
  BUFX3 U233 ( .A(P13[7]), .Y(P12[5]) );
  XOR2X1 U234 ( .A(n59), .B(n60), .Y(P15[1]) );
  BUFX3 U235 ( .A(P1[5]), .Y(P3[9]) );
  XNOR2X1 U236 ( .A(n19), .B(n33), .Y(P7[1]) );
  XOR2X1 U237 ( .A(n84), .B(n90), .Y(P10[1]) );
  XNOR2X1 U238 ( .A(n19), .B(P4[3]), .Y(P9[2]) );
  XNOR2X1 U239 ( .A(n38), .B(P7[3]), .Y(P12[2]) );
  XNOR2XL U240 ( .A(n66), .B(n67), .Y(P14[2]) );
  XNOR2X1 U241 ( .A(n73), .B(n49), .Y(P13[2]) );
  XOR2X1 U242 ( .A(n52), .B(n69), .Y(P11[3]) );
  XOR2X1 U243 ( .A(n51), .B(n58), .Y(P14[1]) );
  BUFX3 U244 ( .A(P10[12]), .Y(P6[4]) );
  BUFX3 U245 ( .A(P10[12]), .Y(P8[8]) );
  BUFX3 U246 ( .A(P10[12]), .Y(P7[6]) );
  BUFX3 U247 ( .A(P12[12]), .Y(P11[10]) );
  BUFX3 U248 ( .A(P12[12]), .Y(P10[8]) );
  BUFX3 U249 ( .A(P12[12]), .Y(P9[6]) );
  BUFX3 U250 ( .A(P12[12]), .Y(P8[4]) );
  BUFX3 U251 ( .A(P1[4]), .Y(P3[8]) );
  BUFX3 U252 ( .A(P1[4]), .Y(P2[6]) );
  BUFX3 U253 ( .A(P5[10]), .Y(P3[6]) );
  BUFX3 U254 ( .A(P13[7]), .Y(P15[11]) );
  BUFX3 U255 ( .A(P15[0]), .Y(P14[11]) );
  BUFX3 U256 ( .A(P15[0]), .Y(P11[5]) );
  BUFX3 U257 ( .A(P15[0]), .Y(P13[9]) );
  BUFX3 U258 ( .A(P15[0]), .Y(P12[7]) );
  BUFX3 U259 ( .A(P13[7]), .Y(P14[9]) );
  BUFX3 U260 ( .A(P13[10]), .Y(P12[8]) );
  BUFX3 U261 ( .A(P13[10]), .Y(P11[6]) );
  BUFX3 U262 ( .A(P13[10]), .Y(P10[4]) );
  BUFX3 U263 ( .A(P13[10]), .Y(P14[12]) );
  XNOR2XL U264 ( .A(n35), .B(P2[10]), .Y(n51) );
  CLKBUFXL U265 ( .A(P2[10]), .Y(P3[12]) );
  INVX1 U266 ( .A(n53), .Y(P2[11]) );
  CLKBUFXL U267 ( .A(P2[10]), .Y(P1[8]) );
  XOR2X1 U268 ( .A(n15), .B(n16), .Y(P9[4]) );
  XNOR2X1 U269 ( .A(n17), .B(b[10]), .Y(n16) );
  XNOR2X1 U270 ( .A(b[11]), .B(b[8]), .Y(n89) );
  XNOR2X1 U271 ( .A(b[2]), .B(n28), .Y(n36) );
  INVX1 U272 ( .A(b[11]), .Y(n35) );
  XNOR2X1 U273 ( .A(b[2]), .B(n38), .Y(n59) );
  XNOR2X1 U274 ( .A(n83), .B(n84), .Y(n52) );
  XNOR2X1 U275 ( .A(n32), .B(P1[3]), .Y(n26) );
  INVX1 U276 ( .A(b[0]), .Y(n42) );
  XNOR2XL U277 ( .A(b[11]), .B(n19), .Y(P2[2]) );
  XOR2X1 U278 ( .A(n21), .B(b[6]), .Y(n6) );
  BUFX3 U279 ( .A(b[5]), .Y(P2[9]) );
  XOR2X1 U280 ( .A(n18), .B(n36), .Y(P10[3]) );
  XNOR2XL U281 ( .A(b[1]), .B(n56), .Y(P15[3]) );
  BUFX3 U282 ( .A(b[3]), .Y(n205) );
  CLKBUFXL U283 ( .A(b[9]), .Y(P2[0]) );
  BUFX3 U284 ( .A(b[8]), .Y(P2[12]) );
  CLKBUFXL U285 ( .A(b[9]), .Y(P1[11]) );
  XNOR2X1 U286 ( .A(n38), .B(b[11]), .Y(n90) );
  CLKBUFXL U287 ( .A(b[10]), .Y(P1[12]) );
  BUFX3 U288 ( .A(b[8]), .Y(P1[10]) );
endmodule


module multiplier_column1_p16 ( b, P1, P2, P3, P4, P5, P6, P7, P8, P9, P10, 
        P11, P12, P13, P14, P15, P16 );
  input [12:0] b;
  output [12:0] P1;
  output [12:0] P2;
  output [12:0] P3;
  output [12:0] P4;
  output [12:0] P5;
  output [12:0] P6;
  output [12:0] P7;
  output [12:0] P8;
  output [12:0] P9;
  output [12:0] P10;
  output [12:0] P11;
  output [12:0] P12;
  output [12:0] P13;
  output [12:0] P14;
  output [12:0] P15;
  output [12:0] P16;
  wire   b_0, P2_1, P3_1, P4_1, P5_1, P6_1, P7_1, P8_1, P9_1, P10_1, P11_1,
         P12_1, P13_1, P14_1, P15_1, P16_1, n6, n7, n8, n9, n11, n12, n13, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n25, n26, n27, n28, n29, n3,
         n33, n34, n35, n36, n37, n154, n194;
  assign b_0 = b[0];
  assign P2[1] = P2_1;
  assign P3[1] = P3_1;
  assign P4[1] = P4_1;
  assign P5[1] = P5_1;
  assign P7[2] = P6_1;
  assign P7[1] = P7_1;
  assign P8[1] = P8_1;
  assign P10[2] = P9_1;
  assign P11[2] = P10_1;
  assign P12[2] = P11_1;
  assign P12[1] = P12_1;
  assign P13[1] = P13_1;
  assign P15[2] = P14_1;
  assign P15[1] = P15_1;
  assign P16[1] = P16_1;

  XOR2X1 U1 ( .A(P2[0]), .B(P1[3]), .Y(P10[12]) );
  XOR2X1 U2 ( .A(P5[10]), .B(P7[3]), .Y(P14[10]) );
  INVX1 U3 ( .A(b[5]), .Y(n3) );
  INVX1 U4 ( .A(n3), .Y(P5[10]) );
  BUFX3 U5 ( .A(n194), .Y(P6[0]) );
  BUFX3 U6 ( .A(n33), .Y(P9[9]) );
  BUFX3 U7 ( .A(n37), .Y(P4[7]) );
  XNOR2XL U8 ( .A(n23), .B(b[12]), .Y(n37) );
  BUFX1 U9 ( .A(P13[7]), .Y(P10[4]) );
  XOR2XL U10 ( .A(P1[5]), .B(n37), .Y(P10_1) );
  CLKBUFXL U11 ( .A(n37), .Y(P1[4]) );
  CLKBUFXL U12 ( .A(n37), .Y(P9[12]) );
  CLKBUFXL U13 ( .A(n37), .Y(P3[6]) );
  CLKBUFXL U14 ( .A(n37), .Y(P2[5]) );
  CLKBUFXL U15 ( .A(P16[0]), .Y(P15[12]) );
  CLKBUFXL U16 ( .A(P16[0]), .Y(P7[4]) );
  CLKBUFXL U17 ( .A(P16[0]), .Y(P9[6]) );
  CLKBUFXL U18 ( .A(P16[0]), .Y(P8[5]) );
  CLKBUFXL U19 ( .A(P16[0]), .Y(P12[9]) );
  CLKBUFXL U20 ( .A(P16[0]), .Y(P10[7]) );
  CLKBUFXL U21 ( .A(P16[0]), .Y(P11[8]) );
  CLKBUFXL U22 ( .A(P9[9]), .Y(P6[6]) );
  CLKBUFXL U23 ( .A(n33), .Y(P8[8]) );
  CLKBUFXL U24 ( .A(P5[4]), .Y(P11[10]) );
  CLKBUFXL U25 ( .A(n33), .Y(P11[11]) );
  BUFX3 U26 ( .A(P3[4]), .Y(P9[10]) );
  XNOR2X1 U27 ( .A(n6), .B(P6[3]), .Y(P16[0]) );
  CLKBUFXL U28 ( .A(n33), .Y(P4[4]) );
  CLKBUFXL U29 ( .A(n33), .Y(P5[5]) );
  CLKBUFXL U30 ( .A(n33), .Y(P7[7]) );
  CLKBUFXL U31 ( .A(P15[0]), .Y(P7[5]) );
  CLKBUFXL U32 ( .A(P15[0]), .Y(P9[7]) );
  CLKBUFXL U33 ( .A(P15[0]), .Y(P11[9]) );
  CLKBUFXL U34 ( .A(P15[0]), .Y(P13[11]) );
  CLKBUFXL U35 ( .A(P15[0]), .Y(P8[6]) );
  CLKBUFXL U36 ( .A(P15[0]), .Y(P12[10]) );
  CLKBUFXL U37 ( .A(P5[4]), .Y(P6[5]) );
  CLKBUFXL U38 ( .A(P5[4]), .Y(P10[9]) );
  CLKBUFXL U39 ( .A(P5[4]), .Y(P7[6]) );
  CLKBUFXL U40 ( .A(P5[4]), .Y(P13[12]) );
  CLKBUFXL U41 ( .A(P5[4]), .Y(P12[11]) );
  XNOR2XL U42 ( .A(n6), .B(P2[2]), .Y(n9) );
  CLKBUFXL U43 ( .A(P2[2]), .Y(P1[1]) );
  CLKBUFXL U44 ( .A(P4_1), .Y(P5[2]) );
  CLKBUFXL U45 ( .A(n33), .Y(P12[12]) );
  CLKBUFXL U46 ( .A(P16[0]), .Y(P13[10]) );
  CLKBUFXL U47 ( .A(n33), .Y(P10[10]) );
  CLKBUFXL U48 ( .A(P2_1), .Y(P3[2]) );
  CLKBUFXL U49 ( .A(P3_1), .Y(P4[2]) );
  XNOR2X1 U50 ( .A(n7), .B(P2[3]), .Y(P3[4]) );
  XOR2X1 U51 ( .A(n194), .B(P5[3]), .Y(P15[0]) );
  XOR2X1 U52 ( .A(P1[9]), .B(P4[3]), .Y(P5[4]) );
  XOR2X1 U53 ( .A(P3[3]), .B(P1[10]), .Y(n33) );
  CLKBUFXL U54 ( .A(P1[10]), .Y(P4[0]) );
  CLKBUFXL U55 ( .A(P1[10]), .Y(P3[12]) );
  CLKBUFXL U56 ( .A(P1[10]), .Y(P2[11]) );
  XOR2XL U57 ( .A(b[2]), .B(b[12]), .Y(P1[3]) );
  XNOR2XL U58 ( .A(P1[9]), .B(n7), .Y(n17) );
  XOR2X1 U59 ( .A(n34), .B(P2[3]), .Y(n21) );
  XOR2X1 U60 ( .A(b_0), .B(P1[10]), .Y(n34) );
  XOR2X1 U61 ( .A(P16_1), .B(n35), .Y(P16[3]) );
  XOR2X1 U62 ( .A(b_0), .B(n194), .Y(n35) );
  XOR2X1 U63 ( .A(n33), .B(n36), .Y(P15[3]) );
  XOR2X1 U64 ( .A(b[1]), .B(P6_1), .Y(n36) );
  XNOR2XL U65 ( .A(n13), .B(P1[10]), .Y(n12) );
  CLKBUFXL U66 ( .A(b[10]), .Y(P2[12]) );
  CLKBUFXL U67 ( .A(b[10]), .Y(P3[0]) );
  CLKBUFXL U68 ( .A(b[10]), .Y(P1[11]) );
  CLKBUFXL U69 ( .A(b[12]), .Y(P1[0]) );
  BUFX3 U70 ( .A(P10[12]), .Y(P9[11]) );
  BUFX3 U71 ( .A(P5[4]), .Y(P8[7]) );
  INVX1 U72 ( .A(n154), .Y(P9[0]) );
  BUFX3 U73 ( .A(P10[12]), .Y(P6[8]) );
  INVX1 U74 ( .A(n154), .Y(P6[10]) );
  BUFX3 U75 ( .A(P3[4]), .Y(P4[5]) );
  XOR2X1 U76 ( .A(P4_1), .B(n8), .Y(n20) );
  BUFX3 U77 ( .A(P12[4]), .Y(P15[7]) );
  INVX1 U78 ( .A(n154), .Y(P7[11]) );
  BUFX3 U79 ( .A(P3[4]), .Y(P6[7]) );
  BUFX3 U80 ( .A(P3[4]), .Y(P12[0]) );
  BUFX3 U81 ( .A(P9[4]), .Y(P11[6]) );
  BUFX3 U82 ( .A(P3[4]), .Y(P11[12]) );
  BUFX3 U83 ( .A(P9[4]), .Y(P10[5]) );
  BUFX3 U84 ( .A(P15[0]), .Y(P10[8]) );
  BUFX3 U85 ( .A(P9_1), .Y(P9[1]) );
  BUFX3 U86 ( .A(P7_1), .Y(P8[2]) );
  INVX1 U87 ( .A(n154), .Y(P4[8]) );
  BUFX3 U88 ( .A(P13[4]), .Y(P14[5]) );
  BUFX3 U89 ( .A(P13[7]), .Y(P15[9]) );
  BUFX3 U90 ( .A(P12[5]), .Y(P14[7]) );
  BUFX3 U91 ( .A(P9[4]), .Y(P15[10]) );
  BUFX3 U92 ( .A(P12[5]), .Y(P11[4]) );
  BUFX3 U93 ( .A(P9[4]), .Y(P12[7]) );
  BUFX3 U94 ( .A(P5[4]), .Y(P14[0]) );
  BUFX3 U95 ( .A(P12[4]), .Y(P13[5]) );
  BUFX3 U96 ( .A(P13[7]), .Y(P14[8]) );
  BUFX3 U97 ( .A(P14[10]), .Y(P11[7]) );
  BUFX3 U98 ( .A(P14[10]), .Y(P8[4]) );
  BUFX3 U99 ( .A(P5[4]), .Y(P9[8]) );
  BUFX3 U100 ( .A(P16[0]), .Y(P14[11]) );
  BUFX3 U101 ( .A(P9[4]), .Y(P13[8]) );
  BUFX3 U102 ( .A(P15[0]), .Y(P14[12]) );
  BUFX3 U103 ( .A(P13[7]), .Y(P12[6]) );
  BUFX3 U104 ( .A(P13[7]), .Y(P11[5]) );
  BUFX3 U105 ( .A(P14[10]), .Y(P12[8]) );
  BUFX3 U106 ( .A(P3[4]), .Y(P10[11]) );
  BUFX3 U107 ( .A(P14[10]), .Y(P15[11]) );
  BUFX3 U108 ( .A(P10[12]), .Y(P11[0]) );
  XOR2X1 U109 ( .A(n27), .B(n28), .Y(P12[3]) );
  BUFX3 U110 ( .A(P10[12]), .Y(P8[10]) );
  INVX1 U111 ( .A(n154), .Y(P2[6]) );
  BUFX3 U112 ( .A(P12_1), .Y(P13[2]) );
  BUFX3 U113 ( .A(P9[9]), .Y(P13[0]) );
  BUFX3 U114 ( .A(P10[12]), .Y(P7[9]) );
  BUFX3 U115 ( .A(P10[12]), .Y(P4[6]) );
  BUFX3 U116 ( .A(P3[4]), .Y(P8[9]) );
  BUFX3 U117 ( .A(P15[0]), .Y(P6[4]) );
  BUFX3 U118 ( .A(P3[4]), .Y(P7[8]) );
  BUFX3 U119 ( .A(P3[4]), .Y(P5[6]) );
  BUFX3 U120 ( .A(P10[12]), .Y(P5[7]) );
  BUFX3 U121 ( .A(P9[4]), .Y(P16[11]) );
  BUFX3 U122 ( .A(P13[7]), .Y(P16[10]) );
  BUFX3 U123 ( .A(P12[5]), .Y(P16[9]) );
  BUFX3 U124 ( .A(P9[4]), .Y(P14[9]) );
  BUFX3 U125 ( .A(P12[4]), .Y(P16[8]) );
  BUFX3 U126 ( .A(P12[5]), .Y(P15[8]) );
  BUFX3 U127 ( .A(P12[5]), .Y(P13[6]) );
  BUFX3 U128 ( .A(P13[4]), .Y(P16[7]) );
  BUFX3 U129 ( .A(P12[4]), .Y(P14[6]) );
  BUFX3 U130 ( .A(P13[4]), .Y(P15[6]) );
  INVX1 U131 ( .A(n154), .Y(P3[7]) );
  BUFX3 U132 ( .A(P14[10]), .Y(P16[12]) );
  BUFX3 U133 ( .A(P14_1), .Y(P14[1]) );
  BUFX3 U134 ( .A(P10_1), .Y(P10[1]) );
  BUFX3 U135 ( .A(P14[10]), .Y(P10[6]) );
  BUFX3 U136 ( .A(P14[10]), .Y(P9[5]) );
  BUFX3 U137 ( .A(P14[10]), .Y(P13[9]) );
  BUFX3 U138 ( .A(P10[12]), .Y(P3[5]) );
  BUFX3 U139 ( .A(P5_1), .Y(P6[2]) );
  INVX1 U140 ( .A(n154), .Y(P5[9]) );
  XOR2X1 U141 ( .A(P1[5]), .B(P8[3]), .Y(P9[4]) );
  XOR2X1 U142 ( .A(P9[3]), .B(n37), .Y(P13[7]) );
  XOR2X1 U143 ( .A(n19), .B(n29), .Y(P12[5]) );
  XOR2X1 U144 ( .A(n25), .B(n26), .Y(P12[4]) );
  XOR2X1 U145 ( .A(n21), .B(n22), .Y(P13[4]) );
  XNOR2X1 U146 ( .A(n23), .B(P1[5]), .Y(n22) );
  XOR2X1 U147 ( .A(n194), .B(P1[9]), .Y(P6_1) );
  XNOR2X1 U148 ( .A(n7), .B(P2[0]), .Y(P3_1) );
  XNOR2X1 U149 ( .A(P1[10]), .B(n7), .Y(P4_1) );
  XNOR2X1 U150 ( .A(n6), .B(n194), .Y(P7_1) );
  XNOR2X1 U151 ( .A(b[5]), .B(n6), .Y(P8_1) );
  XOR2X1 U152 ( .A(P1[10]), .B(P1[9]), .Y(P5_1) );
  XOR2X1 U153 ( .A(P1[9]), .B(P3_1), .Y(P5[3]) );
  XOR2X1 U154 ( .A(n194), .B(P4_1), .Y(P6[3]) );
  XOR2X1 U155 ( .A(b[5]), .B(P1[5]), .Y(P9_1) );
  XOR2X1 U156 ( .A(P3[9]), .B(P5_1), .Y(P7[3]) );
  BUFX3 U157 ( .A(P3[9]), .Y(P5[11]) );
  XOR2X1 U158 ( .A(P7[3]), .B(P2[0]), .Y(P16_1) );
  XNOR2X1 U159 ( .A(n15), .B(P5[3]), .Y(P14_1) );
  XOR2X1 U160 ( .A(P1[3]), .B(n25), .Y(P12_1) );
  XNOR2X1 U161 ( .A(n23), .B(P8_1), .Y(n29) );
  XOR2X1 U162 ( .A(P9_1), .B(P1[3]), .Y(n26) );
  XOR2X1 U163 ( .A(P1[10]), .B(P2_1), .Y(P4[3]) );
  XOR2X1 U164 ( .A(P5[10]), .B(P6_1), .Y(P8[3]) );
  XOR2X1 U165 ( .A(P1[5]), .B(P7_1), .Y(P9[3]) );
  INVX1 U166 ( .A(P3[9]), .Y(n6) );
  BUFX3 U167 ( .A(P5[10]), .Y(P8[0]) );
  BUFX3 U168 ( .A(P3[9]), .Y(P7[0]) );
  BUFX3 U169 ( .A(P5[10]), .Y(P7[12]) );
  BUFX3 U170 ( .A(P3[9]), .Y(P6[12]) );
  BUFX3 U171 ( .A(P6[0]), .Y(P5[12]) );
  BUFX3 U172 ( .A(P3[9]), .Y(P4[10]) );
  BUFX3 U173 ( .A(P6_1), .Y(P6[1]) );
  XOR2X1 U174 ( .A(n8), .B(n9), .Y(P16[4]) );
  XOR2X1 U175 ( .A(P3_1), .B(n37), .Y(n28) );
  BUFX3 U176 ( .A(n194), .Y(P2[9]) );
  XOR2X1 U177 ( .A(n19), .B(n20), .Y(P14[3]) );
  BUFX3 U178 ( .A(P4[7]), .Y(P10[0]) );
  INVX1 U179 ( .A(n154), .Y(P8[12]) );
  XOR2X1 U180 ( .A(P2[0]), .B(n26), .Y(P11[3]) );
  BUFX3 U181 ( .A(P4[7]), .Y(P7[10]) );
  BUFX3 U182 ( .A(P5[10]), .Y(P6[11]) );
  BUFX3 U183 ( .A(P1[9]), .Y(P5[0]) );
  BUFX3 U184 ( .A(P5[10]), .Y(P4[9]) );
  BUFX3 U185 ( .A(n194), .Y(P4[11]) );
  BUFX3 U186 ( .A(P5[10]), .Y(P3[8]) );
  BUFX3 U187 ( .A(P10[12]), .Y(P2[4]) );
  BUFX3 U188 ( .A(P5[10]), .Y(P2[7]) );
  BUFX3 U189 ( .A(P3[9]), .Y(P2[8]) );
  XOR2X1 U190 ( .A(n33), .B(P11_1), .Y(P13[3]) );
  BUFX3 U191 ( .A(P4[7]), .Y(P5[8]) );
  BUFX3 U192 ( .A(P8_1), .Y(P9[2]) );
  BUFX3 U193 ( .A(P11_1), .Y(P11[1]) );
  BUFX3 U194 ( .A(P15_1), .Y(P16[2]) );
  BUFX3 U195 ( .A(P13_1), .Y(P14[2]) );
  XNOR2X1 U196 ( .A(n13), .B(P1[9]), .Y(n8) );
  BUFX3 U197 ( .A(P1[9]), .Y(P4[12]) );
  BUFX3 U198 ( .A(P1[9]), .Y(P2[10]) );
  XNOR2X1 U199 ( .A(P1[5]), .B(n13), .Y(n27) );
  INVX1 U200 ( .A(P1[5]), .Y(n154) );
  BUFX3 U201 ( .A(P14[4]), .Y(P16[6]) );
  BUFX3 U202 ( .A(P14[4]), .Y(P15[5]) );
  BUFX3 U203 ( .A(P16[5]), .Y(P15[4]) );
  CLKBUFXL U204 ( .A(n37), .Y(P8[11]) );
  CLKBUFXL U205 ( .A(n37), .Y(P6[9]) );
  BUFX3 U206 ( .A(P1[9]), .Y(P3[11]) );
  BUFX3 U207 ( .A(n194), .Y(P3[10]) );
  BUFX3 U208 ( .A(P5[10]), .Y(P1[6]) );
  BUFX3 U209 ( .A(P6[0]), .Y(P1[8]) );
  BUFX3 U210 ( .A(P3[9]), .Y(P1[7]) );
  XNOR2X1 U211 ( .A(n15), .B(b[12]), .Y(P2[2]) );
  XOR2X1 U212 ( .A(b[12]), .B(P2[0]), .Y(P2_1) );
  XOR2X1 U213 ( .A(P2[0]), .B(b[1]), .Y(P2[3]) );
  XOR2X1 U214 ( .A(b[2]), .B(P2[0]), .Y(n19) );
  XOR2X1 U215 ( .A(b[12]), .B(P6[3]), .Y(P15_1) );
  XOR2X1 U216 ( .A(b[12]), .B(n21), .Y(P13_1) );
  INVX1 U217 ( .A(b[10]), .Y(n7) );
  XOR2X1 U218 ( .A(b[10]), .B(P2[2]), .Y(P3[3]) );
  XNOR2X1 U219 ( .A(n7), .B(b[1]), .Y(n25) );
  BUFX3 U220 ( .A(b[7]), .Y(n194) );
  BUFX3 U221 ( .A(b[8]), .Y(P1[9]) );
  BUFX3 U222 ( .A(b[6]), .Y(P3[9]) );
  XOR2X1 U223 ( .A(b[12]), .B(n29), .Y(P10[3]) );
  BUFX3 U224 ( .A(b[9]), .Y(P1[10]) );
  BUFX3 U225 ( .A(b[11]), .Y(P2[0]) );
  INVX1 U226 ( .A(b[3]), .Y(n23) );
  INVX1 U227 ( .A(b_0), .Y(n15) );
  BUFX3 U228 ( .A(b[4]), .Y(P1[5]) );
  XOR2X1 U229 ( .A(n16), .B(n17), .Y(P14[4]) );
  XOR2X1 U230 ( .A(b[2]), .B(n18), .Y(n16) );
  XNOR2X1 U231 ( .A(n15), .B(b[3]), .Y(n18) );
  XOR2X1 U232 ( .A(b[3]), .B(n19), .Y(P11_1) );
  XOR2X1 U233 ( .A(n11), .B(n12), .Y(P16[5]) );
  XOR2X1 U234 ( .A(b[2]), .B(n194), .Y(n11) );
  INVX1 U235 ( .A(b[1]), .Y(n13) );
  BUFX3 U236 ( .A(b[1]), .Y(P1[2]) );
  BUFX3 U237 ( .A(P2[0]), .Y(P1[12]) );
endmodule


module mux13_13_8 ( a, b, sel, enable, out, clk, reset );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel, enable, clk, reset;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N83,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29;

  EDFFX1 \out_reg[12]  ( .D(N29), .E(N83), .CK(clk), .Q(out[12]) );
  EDFFX1 \out_reg[11]  ( .D(N28), .E(N83), .CK(clk), .Q(out[11]) );
  EDFFX1 \out_reg[10]  ( .D(N27), .E(N83), .CK(clk), .Q(out[10]) );
  EDFFX1 \out_reg[9]  ( .D(N26), .E(N83), .CK(clk), .Q(out[9]) );
  EDFFX1 \out_reg[8]  ( .D(N25), .E(N83), .CK(clk), .Q(out[8]) );
  EDFFX1 \out_reg[7]  ( .D(N24), .E(N83), .CK(clk), .Q(out[7]) );
  EDFFX1 \out_reg[6]  ( .D(N23), .E(N83), .CK(clk), .Q(out[6]) );
  EDFFX1 \out_reg[5]  ( .D(N22), .E(N83), .CK(clk), .Q(out[5]) );
  EDFFX1 \out_reg[4]  ( .D(N21), .E(N83), .CK(clk), .Q(out[4]) );
  EDFFX1 \out_reg[3]  ( .D(N20), .E(N83), .CK(clk), .Q(out[3]) );
  EDFFX1 \out_reg[2]  ( .D(N19), .E(N83), .CK(clk), .Q(out[2]) );
  EDFFX1 \out_reg[1]  ( .D(N18), .E(N83), .CK(clk), .Q(out[1]) );
  EDFFX1 \out_reg[0]  ( .D(N17), .E(N83), .CK(clk), .Q(out[0]) );
  NAND2BX1 U3 ( .AN(enable), .B(reset), .Y(N83) );
  NOR2BX1 U4 ( .AN(reset), .B(sel), .Y(n16) );
  AND2X2 U5 ( .A(sel), .B(reset), .Y(n17) );
  INVX1 U6 ( .A(n29), .Y(N17) );
  AOI22X1 U7 ( .A0(b[0]), .A1(n16), .B0(a[0]), .B1(n17), .Y(n29) );
  INVX1 U8 ( .A(n28), .Y(N18) );
  AOI22X1 U9 ( .A0(b[1]), .A1(n16), .B0(a[1]), .B1(n17), .Y(n28) );
  INVX1 U10 ( .A(n27), .Y(N19) );
  AOI22X1 U11 ( .A0(b[2]), .A1(n16), .B0(a[2]), .B1(n17), .Y(n27) );
  INVX1 U12 ( .A(n26), .Y(N20) );
  AOI22X1 U13 ( .A0(b[3]), .A1(n16), .B0(a[3]), .B1(n17), .Y(n26) );
  INVX1 U14 ( .A(n25), .Y(N21) );
  AOI22X1 U15 ( .A0(b[4]), .A1(n16), .B0(a[4]), .B1(n17), .Y(n25) );
  INVX1 U16 ( .A(n24), .Y(N22) );
  AOI22X1 U17 ( .A0(b[5]), .A1(n16), .B0(a[5]), .B1(n17), .Y(n24) );
  INVX1 U18 ( .A(n23), .Y(N23) );
  AOI22X1 U19 ( .A0(b[6]), .A1(n16), .B0(a[6]), .B1(n17), .Y(n23) );
  INVX1 U20 ( .A(n22), .Y(N24) );
  AOI22X1 U21 ( .A0(b[7]), .A1(n16), .B0(a[7]), .B1(n17), .Y(n22) );
  INVX1 U22 ( .A(n21), .Y(N25) );
  AOI22X1 U23 ( .A0(b[8]), .A1(n16), .B0(a[8]), .B1(n17), .Y(n21) );
  INVX1 U24 ( .A(n20), .Y(N26) );
  AOI22X1 U25 ( .A0(b[9]), .A1(n16), .B0(a[9]), .B1(n17), .Y(n20) );
  INVX1 U26 ( .A(n19), .Y(N27) );
  AOI22X1 U27 ( .A0(b[10]), .A1(n16), .B0(a[10]), .B1(n17), .Y(n19) );
  INVX1 U28 ( .A(n18), .Y(N28) );
  AOI22X1 U29 ( .A0(b[11]), .A1(n16), .B0(a[11]), .B1(n17), .Y(n18) );
  INVX1 U30 ( .A(n15), .Y(N29) );
  AOI22X1 U31 ( .A0(b[12]), .A1(n16), .B0(a[12]), .B1(n17), .Y(n15) );
endmodule


module multiply_7163 ( a, c );
  input [12:0] a;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;

  XOR2X1 U1 ( .A(n1), .B(n2), .Y(c[9]) );
  XNOR2X1 U2 ( .A(n3), .B(n4), .Y(n2) );
  XOR2X1 U3 ( .A(n17), .B(n14), .Y(c[11]) );
  XNOR2X1 U4 ( .A(n6), .B(n4), .Y(n14) );
  XOR2X1 U5 ( .A(n4), .B(n11), .Y(n5) );
  XNOR2X1 U6 ( .A(n3), .B(n17), .Y(n8) );
  XNOR2X1 U7 ( .A(n6), .B(n11), .Y(n24) );
  XNOR2X1 U8 ( .A(n3), .B(n5), .Y(n21) );
  XOR2X1 U9 ( .A(n1), .B(n11), .Y(n10) );
  XOR2X1 U10 ( .A(n22), .B(n23), .Y(c[1]) );
  XOR2X1 U11 ( .A(a[9]), .B(a[6]), .Y(n22) );
  XOR2X1 U12 ( .A(a[6]), .B(n5), .Y(c[8]) );
  XOR2X1 U13 ( .A(n17), .B(n26), .Y(c[10]) );
  XOR2X1 U14 ( .A(a[6]), .B(n1), .Y(n26) );
  XOR2X1 U15 ( .A(n8), .B(n27), .Y(c[0]) );
  XOR2X1 U16 ( .A(a[1]), .B(n11), .Y(n27) );
  XOR2X1 U17 ( .A(n15), .B(n16), .Y(c[3]) );
  XOR2X1 U18 ( .A(a[4]), .B(n19), .Y(n15) );
  XOR2X1 U19 ( .A(n12), .B(n13), .Y(c[4]) );
  XOR2X1 U20 ( .A(a[2]), .B(a[12]), .Y(n12) );
  XOR2X1 U21 ( .A(n9), .B(n10), .Y(c[5]) );
  XOR2X1 U22 ( .A(a[3]), .B(a[12]), .Y(n9) );
  XOR2X1 U23 ( .A(a[4]), .B(n8), .Y(c[6]) );
  XNOR2X1 U24 ( .A(n6), .B(n7), .Y(c[7]) );
  XOR2X1 U25 ( .A(a[6]), .B(a[5]), .Y(n7) );
  XOR2X1 U26 ( .A(a[11]), .B(a[4]), .Y(n11) );
  XOR2X1 U27 ( .A(a[1]), .B(a[8]), .Y(n1) );
  XOR2X1 U28 ( .A(a[2]), .B(a[9]), .Y(n17) );
  XOR2X1 U29 ( .A(a[0]), .B(a[7]), .Y(n4) );
  XNOR2X1 U30 ( .A(a[12]), .B(a[5]), .Y(n3) );
  XNOR2X1 U31 ( .A(a[10]), .B(a[3]), .Y(n6) );
  XOR2X1 U32 ( .A(a[1]), .B(n24), .Y(n23) );
  XOR2X1 U33 ( .A(a[8]), .B(a[6]), .Y(n19) );
  XOR2X1 U34 ( .A(a[11]), .B(n14), .Y(n13) );
  XOR2X1 U35 ( .A(n17), .B(n18), .Y(n16) );
  XOR2X1 U36 ( .A(a[3]), .B(a[0]), .Y(n18) );
  XOR2X1 U37 ( .A(n20), .B(n21), .Y(c[2]) );
  XOR2X1 U38 ( .A(a[2]), .B(a[10]), .Y(n20) );
  XOR2X1 U39 ( .A(n24), .B(n25), .Y(c[12]) );
  XOR2X1 U40 ( .A(a[0]), .B(n1), .Y(n25) );
endmodule


module multiply_3196 ( a, c );
  input [12:0] a;
  output [12:0] c;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR2X1 U1 ( .A(n39), .B(n40), .Y(c[0]) );
  XNOR2X1 U2 ( .A(n16), .B(n38), .Y(n40) );
  XOR2X1 U3 ( .A(n19), .B(n31), .Y(c[12]) );
  XNOR2X1 U4 ( .A(n30), .B(n13), .Y(n31) );
  XNOR2X1 U5 ( .A(n16), .B(n5), .Y(n23) );
  XNOR2X1 U6 ( .A(n30), .B(n12), .Y(n4) );
  XNOR2X1 U7 ( .A(n30), .B(n9), .Y(n20) );
  XOR2X1 U8 ( .A(n12), .B(n5), .Y(n8) );
  XNOR2X1 U9 ( .A(n4), .B(n16), .Y(n15) );
  XOR2X1 U10 ( .A(n9), .B(n23), .Y(n22) );
  XOR2X1 U11 ( .A(n23), .B(n38), .Y(n37) );
  XOR2XL U12 ( .A(n12), .B(n13), .Y(n11) );
  XOR2X1 U13 ( .A(n4), .B(n5), .Y(n3) );
  XOR2X1 U14 ( .A(n19), .B(n20), .Y(n18) );
  XOR2X1 U15 ( .A(n20), .B(n24), .Y(n35) );
  XOR2X1 U16 ( .A(n8), .B(n9), .Y(n7) );
  XNOR2X1 U17 ( .A(a[11]), .B(a[4]), .Y(n16) );
  XOR2X1 U18 ( .A(n32), .B(n16), .Y(n13) );
  XOR2X1 U19 ( .A(n33), .B(a[1]), .Y(n32) );
  INVX1 U20 ( .A(a[12]), .Y(n33) );
  XOR2X1 U21 ( .A(n28), .B(n29), .Y(c[1]) );
  XOR2X1 U22 ( .A(n10), .B(n11), .Y(c[7]) );
  XOR2X1 U23 ( .A(a[8]), .B(a[5]), .Y(n10) );
  XOR2X1 U24 ( .A(n34), .B(n35), .Y(c[11]) );
  XOR2X1 U25 ( .A(a[12]), .B(n5), .Y(n34) );
  XOR2X1 U26 ( .A(n14), .B(n15), .Y(c[6]) );
  XOR2X1 U27 ( .A(a[5]), .B(a[0]), .Y(n14) );
  XOR2X1 U28 ( .A(n2), .B(n3), .Y(c[9]) );
  XOR2X1 U29 ( .A(a[1]), .B(a[0]), .Y(n2) );
  XOR2X1 U30 ( .A(n26), .B(n27), .Y(c[2]) );
  XOR2X1 U31 ( .A(a[7]), .B(a[5]), .Y(n26) );
  XOR2X1 U32 ( .A(n21), .B(n22), .Y(c[4]) );
  XOR2X1 U33 ( .A(a[3]), .B(a[1]), .Y(n21) );
  XOR2X1 U34 ( .A(n17), .B(n18), .Y(c[5]) );
  XOR2X1 U35 ( .A(a[4]), .B(a[12]), .Y(n17) );
  XOR2X1 U36 ( .A(n6), .B(n7), .Y(c[8]) );
  XOR2X1 U37 ( .A(a[12]), .B(a[0]), .Y(n6) );
  XOR2X1 U38 ( .A(n36), .B(n37), .Y(c[10]) );
  XOR2X1 U39 ( .A(a[2]), .B(a[1]), .Y(n36) );
  XOR2X1 U40 ( .A(a[8]), .B(a[9]), .Y(n5) );
  XOR2X1 U41 ( .A(a[2]), .B(a[5]), .Y(n9) );
  XOR2X1 U42 ( .A(a[6]), .B(a[7]), .Y(n12) );
  XOR2X1 U43 ( .A(a[10]), .B(a[7]), .Y(n38) );
  XNOR2X1 U44 ( .A(a[10]), .B(a[3]), .Y(n30) );
  XOR2X1 U45 ( .A(a[11]), .B(a[0]), .Y(n24) );
  XOR2X1 U46 ( .A(a[6]), .B(a[9]), .Y(n19) );
  XOR2X1 U47 ( .A(a[2]), .B(n4), .Y(n29) );
  XOR2X1 U48 ( .A(a[3]), .B(n23), .Y(n27) );
  XOR2X1 U49 ( .A(a[12]), .B(n9), .Y(n39) );
  XOR2X1 U50 ( .A(a[8]), .B(a[4]), .Y(n28) );
  XOR2X1 U51 ( .A(n24), .B(n25), .Y(c[3]) );
  XOR2X1 U52 ( .A(a[2]), .B(n8), .Y(n25) );
endmodule


module multiply_7420 ( a, c );
  input [12:0] a;
  output [12:0] c;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;

  XOR2X1 U1 ( .A(n25), .B(n4), .Y(n22) );
  XOR2X1 U2 ( .A(n21), .B(n22), .Y(n20) );
  XNOR2X1 U3 ( .A(n32), .B(n21), .Y(n6) );
  XNOR2X1 U4 ( .A(n30), .B(n25), .Y(n9) );
  XOR2X1 U5 ( .A(n5), .B(n9), .Y(n27) );
  XNOR2X1 U6 ( .A(n32), .B(n4), .Y(n13) );
  XNOR2X1 U7 ( .A(n25), .B(n6), .Y(n17) );
  XOR2X1 U8 ( .A(n5), .B(n29), .Y(n16) );
  XNOR2X1 U9 ( .A(n30), .B(n21), .Y(n29) );
  XOR2X1 U10 ( .A(n6), .B(n5), .Y(n12) );
  XOR2X1 U11 ( .A(n4), .B(n9), .Y(n8) );
  XOR2X1 U12 ( .A(n15), .B(n35), .Y(c[0]) );
  XNOR2X1 U13 ( .A(n30), .B(n13), .Y(n35) );
  XOR2X1 U14 ( .A(n15), .B(n16), .Y(c[5]) );
  XOR2X1 U15 ( .A(n2), .B(n3), .Y(c[9]) );
  XOR2X1 U16 ( .A(n4), .B(n5), .Y(n3) );
  XOR2X1 U17 ( .A(a[5]), .B(a[12]), .Y(n4) );
  XOR2X1 U18 ( .A(n19), .B(n20), .Y(c[3]) );
  XOR2X1 U19 ( .A(a[3]), .B(a[11]), .Y(n19) );
  XOR2X1 U20 ( .A(a[11]), .B(a[6]), .Y(n5) );
  XOR2X1 U21 ( .A(a[1]), .B(a[8]), .Y(n21) );
  XOR2X1 U22 ( .A(a[0]), .B(a[7]), .Y(n25) );
  XOR2X1 U23 ( .A(a[2]), .B(n24), .Y(n30) );
  XOR2X1 U24 ( .A(a[7]), .B(a[4]), .Y(n15) );
  XNOR2X1 U25 ( .A(a[10]), .B(a[3]), .Y(n32) );
  XOR2X1 U26 ( .A(a[4]), .B(a[11]), .Y(n10) );
  XOR2X1 U27 ( .A(a[4]), .B(a[1]), .Y(n34) );
  XOR2X1 U28 ( .A(n22), .B(n31), .Y(c[11]) );
  XOR2X1 U29 ( .A(a[2]), .B(n6), .Y(n31) );
  INVX1 U30 ( .A(a[9]), .Y(n24) );
  XOR2X1 U31 ( .A(n17), .B(n18), .Y(c[4]) );
  XNOR2X1 U32 ( .A(a[5]), .B(a[6]), .Y(n18) );
  XOR2X1 U33 ( .A(a[0]), .B(n6), .Y(n2) );
  XOR2X1 U34 ( .A(n26), .B(n27), .Y(c[1]) );
  XOR2X1 U35 ( .A(a[8]), .B(a[12]), .Y(n26) );
  XOR2X1 U36 ( .A(n17), .B(n23), .Y(c[2]) );
  XOR2X1 U37 ( .A(n24), .B(a[12]), .Y(n23) );
  XOR2X1 U38 ( .A(n13), .B(n14), .Y(c[6]) );
  XOR2X1 U39 ( .A(a[8]), .B(n9), .Y(n14) );
  XOR2X1 U40 ( .A(n11), .B(n12), .Y(c[7]) );
  XOR2X1 U41 ( .A(a[9]), .B(a[4]), .Y(n11) );
  XOR2X1 U42 ( .A(n7), .B(n8), .Y(c[8]) );
  XOR2X1 U43 ( .A(a[10]), .B(n10), .Y(n7) );
  XOR2X1 U44 ( .A(n33), .B(n27), .Y(c[10]) );
  XOR2X1 U45 ( .A(a[12]), .B(n34), .Y(n33) );
  XOR2X1 U46 ( .A(n28), .B(n16), .Y(c[12]) );
  XOR2X1 U47 ( .A(a[4]), .B(a[3]), .Y(n28) );
endmodule


module multiply_3453 ( a, c );
  input [12:0] a;
  output [12:0] c;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34;

  XOR2X1 U1 ( .A(n7), .B(n8), .Y(c[7]) );
  XNOR2X1 U2 ( .A(n12), .B(n5), .Y(n20) );
  XOR2X1 U3 ( .A(n22), .B(n11), .Y(n8) );
  XOR2X1 U4 ( .A(n2), .B(n11), .Y(n25) );
  XNOR2X1 U5 ( .A(n11), .B(n12), .Y(n10) );
  XOR2X1 U6 ( .A(n7), .B(n25), .Y(n24) );
  INVX1 U7 ( .A(n18), .Y(n2) );
  XOR2X1 U8 ( .A(n2), .B(n3), .Y(c[9]) );
  XOR2X1 U9 ( .A(n4), .B(n5), .Y(n3) );
  XOR2X1 U10 ( .A(n22), .B(n31), .Y(c[12]) );
  XOR2X1 U11 ( .A(a[7]), .B(n17), .Y(n31) );
  XOR2X1 U12 ( .A(n17), .B(n34), .Y(c[0]) );
  XOR2X1 U13 ( .A(a[8]), .B(n4), .Y(n34) );
  XOR2X1 U14 ( .A(n23), .B(n24), .Y(c[3]) );
  XOR2X1 U15 ( .A(a[1]), .B(n26), .Y(n23) );
  XOR2X1 U16 ( .A(n8), .B(n32), .Y(c[11]) );
  XOR2X1 U17 ( .A(a[6]), .B(a[1]), .Y(n32) );
  XOR2X1 U18 ( .A(a[10]), .B(a[3]), .Y(n17) );
  XOR2X1 U19 ( .A(a[12]), .B(a[8]), .Y(n11) );
  XOR2X1 U20 ( .A(n11), .B(n29), .Y(c[1]) );
  XOR2X1 U21 ( .A(a[0]), .B(n6), .Y(n29) );
  XOR2X1 U22 ( .A(n20), .B(n21), .Y(c[4]) );
  XOR2X1 U23 ( .A(a[5]), .B(n22), .Y(n21) );
  XOR2X1 U24 ( .A(n9), .B(n10), .Y(c[6]) );
  XOR2X1 U25 ( .A(a[3]), .B(n13), .Y(n9) );
  XNOR2X1 U26 ( .A(a[11]), .B(a[1]), .Y(n12) );
  XOR2X1 U27 ( .A(a[2]), .B(a[9]), .Y(n22) );
  XNOR2X1 U28 ( .A(n30), .B(n17), .Y(n6) );
  XNOR2X1 U29 ( .A(a[9]), .B(a[5]), .Y(n30) );
  XOR2X1 U30 ( .A(a[10]), .B(a[6]), .Y(n5) );
  XNOR2X1 U31 ( .A(a[0]), .B(a[7]), .Y(n18) );
  XOR2X1 U32 ( .A(a[11]), .B(a[4]), .Y(n4) );
  XOR2X1 U33 ( .A(a[4]), .B(a[5]), .Y(n7) );
  XOR2X1 U34 ( .A(a[6]), .B(a[2]), .Y(n19) );
  XOR2X1 U35 ( .A(a[3]), .B(a[2]), .Y(n26) );
  XOR2X1 U36 ( .A(a[7]), .B(a[4]), .Y(n13) );
  XOR2X1 U37 ( .A(a[0]), .B(n20), .Y(n28) );
  XOR2X1 U38 ( .A(n16), .B(n17), .Y(n15) );
  XOR2X1 U39 ( .A(a[11]), .B(n18), .Y(n16) );
  XOR2X1 U40 ( .A(n14), .B(n15), .Y(c[5]) );
  XNOR2X1 U41 ( .A(a[12]), .B(n19), .Y(n14) );
  XOR2X1 U42 ( .A(n27), .B(n28), .Y(c[2]) );
  XOR2X1 U43 ( .A(a[9]), .B(a[4]), .Y(n27) );
  XOR2X1 U44 ( .A(a[6]), .B(n6), .Y(c[8]) );
  XOR2X1 U45 ( .A(n25), .B(n33), .Y(c[10]) );
  XNOR2X1 U46 ( .A(a[5]), .B(n12), .Y(n33) );
endmodule


module multiply_7677 ( a, c );
  input [12:0] a;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;

  XNOR2X1 U1 ( .A(n10), .B(n8), .Y(n15) );
  XOR2X1 U2 ( .A(n15), .B(n18), .Y(n17) );
  XOR2X1 U3 ( .A(n3), .B(n21), .Y(n20) );
  XOR2X1 U4 ( .A(n19), .B(n20), .Y(c[1]) );
  XOR2X1 U5 ( .A(n1), .B(n22), .Y(n19) );
  XOR2X1 U6 ( .A(n12), .B(n15), .Y(c[3]) );
  XOR2X1 U7 ( .A(a[8]), .B(n21), .Y(c[11]) );
  XOR2X1 U8 ( .A(n16), .B(n17), .Y(c[2]) );
  XOR2X1 U9 ( .A(n3), .B(n25), .Y(c[0]) );
  XOR2X1 U10 ( .A(a[6]), .B(a[4]), .Y(n25) );
  XNOR2X1 U11 ( .A(n10), .B(n24), .Y(c[10]) );
  XOR2X1 U12 ( .A(a[3]), .B(a[1]), .Y(n24) );
  XOR2X1 U13 ( .A(n18), .B(n23), .Y(c[12]) );
  XOR2X1 U14 ( .A(a[9]), .B(a[3]), .Y(n23) );
  XOR2X1 U15 ( .A(a[11]), .B(a[6]), .Y(n1) );
  XOR2X1 U16 ( .A(a[4]), .B(a[2]), .Y(n21) );
  XOR2X1 U17 ( .A(a[10]), .B(a[1]), .Y(n3) );
  XNOR2X1 U18 ( .A(a[12]), .B(a[7]), .Y(n10) );
  XOR2X1 U19 ( .A(a[0]), .B(a[5]), .Y(n18) );
  XOR2X1 U20 ( .A(a[10]), .B(a[9]), .Y(n12) );
  XOR2X1 U21 ( .A(a[3]), .B(a[8]), .Y(n8) );
  XOR2X1 U22 ( .A(a[12]), .B(n7), .Y(n5) );
  XOR2X1 U23 ( .A(a[9]), .B(a[4]), .Y(n7) );
  XOR2X1 U24 ( .A(a[1]), .B(n1), .Y(n14) );
  XOR2X1 U25 ( .A(a[7]), .B(a[5]), .Y(n22) );
  XOR2X1 U26 ( .A(a[2]), .B(n1), .Y(n16) );
  XOR2X1 U27 ( .A(n13), .B(n14), .Y(c[4]) );
  XOR2X1 U28 ( .A(a[9]), .B(a[8]), .Y(n13) );
  XNOR2X1 U29 ( .A(n10), .B(n11), .Y(c[5]) );
  XOR2X1 U30 ( .A(a[2]), .B(n12), .Y(n11) );
  XOR2X1 U31 ( .A(n8), .B(n9), .Y(c[6]) );
  XOR2X1 U32 ( .A(a[11]), .B(a[10]), .Y(n9) );
  XOR2X1 U33 ( .A(n5), .B(n6), .Y(c[7]) );
  XOR2X1 U34 ( .A(a[11]), .B(a[0]), .Y(n6) );
  XOR2X1 U35 ( .A(n3), .B(n4), .Y(c[8]) );
  XOR2X1 U36 ( .A(a[5]), .B(a[12]), .Y(n4) );
  XOR2X1 U37 ( .A(n1), .B(n2), .Y(c[9]) );
  XOR2X1 U38 ( .A(a[2]), .B(a[0]), .Y(n2) );
endmodule


module multiply_3710 ( a, c );
  input [12:0] a;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;

  XOR2X1 U1 ( .A(n10), .B(n14), .Y(c[12]) );
  XNOR2X1 U2 ( .A(n13), .B(n18), .Y(n10) );
  XOR2X1 U3 ( .A(n21), .B(n1), .Y(c[10]) );
  XOR2X1 U4 ( .A(n17), .B(n10), .Y(c[11]) );
  XNOR2X1 U5 ( .A(n26), .B(n7), .Y(n17) );
  XNOR2X1 U6 ( .A(n26), .B(n3), .Y(n14) );
  XNOR2X1 U7 ( .A(n13), .B(n4), .Y(n21) );
  XOR2X1 U8 ( .A(n18), .B(n4), .Y(n5) );
  XNOR2X1 U9 ( .A(n13), .B(n14), .Y(n12) );
  XOR2X1 U10 ( .A(n4), .B(n10), .Y(n9) );
  XOR2X1 U11 ( .A(n3), .B(n10), .Y(n28) );
  XOR2X1 U12 ( .A(n7), .B(n3), .Y(n6) );
  XOR2X1 U13 ( .A(n7), .B(n21), .Y(n20) );
  XOR2X1 U14 ( .A(n17), .B(n18), .Y(n16) );
  XOR2X1 U15 ( .A(n1), .B(n2), .Y(c[9]) );
  XOR2X1 U16 ( .A(n3), .B(n4), .Y(n2) );
  XOR2X1 U17 ( .A(n27), .B(n28), .Y(c[0]) );
  XOR2X1 U18 ( .A(a[6]), .B(a[12]), .Y(n27) );
  XOR2X1 U19 ( .A(a[0]), .B(a[6]), .Y(n4) );
  XOR2X1 U20 ( .A(a[11]), .B(a[5]), .Y(n3) );
  XOR2X1 U21 ( .A(a[10]), .B(a[4]), .Y(n18) );
  XNOR2X1 U22 ( .A(a[7]), .B(n13), .Y(c[1]) );
  XOR2X1 U23 ( .A(n18), .B(n25), .Y(c[2]) );
  XOR2X1 U24 ( .A(a[8]), .B(a[0]), .Y(n25) );
  XOR2X1 U25 ( .A(n15), .B(n16), .Y(c[5]) );
  XOR2X1 U26 ( .A(a[3]), .B(a[11]), .Y(n15) );
  XOR2X1 U27 ( .A(n11), .B(n12), .Y(c[6]) );
  XOR2X1 U28 ( .A(a[4]), .B(a[12]), .Y(n11) );
  XNOR2X1 U29 ( .A(a[3]), .B(a[9]), .Y(n13) );
  XOR2X1 U30 ( .A(a[1]), .B(a[7]), .Y(n7) );
  XOR2X1 U31 ( .A(a[12]), .B(n17), .Y(n1) );
  XNOR2X1 U32 ( .A(a[2]), .B(a[8]), .Y(n26) );
  XOR2X1 U33 ( .A(a[12]), .B(n5), .Y(n24) );
  XOR2X1 U34 ( .A(a[2]), .B(a[12]), .Y(n22) );
  XOR2X1 U35 ( .A(n5), .B(n6), .Y(c[8]) );
  XOR2X1 U36 ( .A(n8), .B(n9), .Y(c[7]) );
  XOR2X1 U37 ( .A(a[5]), .B(a[12]), .Y(n8) );
  XOR2X1 U38 ( .A(n23), .B(n24), .Y(c[3]) );
  XOR2X1 U39 ( .A(a[3]), .B(a[1]), .Y(n23) );
  XOR2X1 U40 ( .A(n19), .B(n20), .Y(c[4]) );
  XOR2X1 U41 ( .A(a[10]), .B(n22), .Y(n19) );
endmodule


module multiply_7934 ( a, c );
  input [12:0] a;
  output [12:0] c;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  XOR2X1 U1 ( .A(n10), .B(n14), .Y(c[4]) );
  XOR2X1 U2 ( .A(n2), .B(n15), .Y(n14) );
  XOR2X1 U3 ( .A(n10), .B(n11), .Y(c[5]) );
  XOR2X1 U4 ( .A(n12), .B(n13), .Y(n11) );
  XOR2X1 U5 ( .A(n8), .B(n9), .Y(c[6]) );
  XOR2X1 U6 ( .A(n4), .B(n23), .Y(c[1]) );
  XOR2X1 U7 ( .A(n13), .B(n15), .Y(n9) );
  XOR2X1 U8 ( .A(n12), .B(n18), .Y(n6) );
  XOR2X1 U9 ( .A(n18), .B(n15), .Y(n17) );
  XOR2X1 U10 ( .A(n8), .B(n15), .Y(n26) );
  XOR2X1 U11 ( .A(a[6]), .B(n23), .Y(c[10]) );
  XOR2X1 U12 ( .A(n30), .B(n31), .Y(c[0]) );
  XOR2X1 U13 ( .A(a[9]), .B(a[2]), .Y(n30) );
  XOR2X1 U14 ( .A(n16), .B(n17), .Y(c[3]) );
  XOR2X1 U15 ( .A(a[10]), .B(n19), .Y(n16) );
  XOR2X1 U16 ( .A(n6), .B(n7), .Y(c[7]) );
  XOR2X1 U17 ( .A(a[6]), .B(a[11]), .Y(n7) );
  XOR2X1 U18 ( .A(n4), .B(n5), .Y(c[8]) );
  XOR2X1 U19 ( .A(a[4]), .B(a[2]), .Y(n5) );
  XOR2X1 U20 ( .A(n2), .B(n3), .Y(c[9]) );
  XOR2X1 U21 ( .A(a[9]), .B(a[5]), .Y(n3) );
  XOR2X1 U22 ( .A(n9), .B(n27), .Y(c[11]) );
  XOR2X1 U23 ( .A(a[7]), .B(a[1]), .Y(n27) );
  XOR2X1 U24 ( .A(n25), .B(n26), .Y(c[12]) );
  XOR2X1 U25 ( .A(a[8]), .B(n12), .Y(n25) );
  XOR2X1 U26 ( .A(a[0]), .B(a[11]), .Y(n15) );
  XOR2X1 U27 ( .A(a[10]), .B(a[5]), .Y(n13) );
  XOR2X1 U28 ( .A(a[12]), .B(a[1]), .Y(n12) );
  XOR2X1 U29 ( .A(a[4]), .B(a[9]), .Y(n10) );
  XNOR2X1 U30 ( .A(n28), .B(n10), .Y(n23) );
  XOR2X1 U31 ( .A(n29), .B(a[10]), .Y(n28) );
  INVX1 U32 ( .A(a[0]), .Y(n29) );
  XOR2X1 U33 ( .A(a[3]), .B(a[7]), .Y(n18) );
  XOR2X1 U34 ( .A(a[2]), .B(a[6]), .Y(n8) );
  XOR2X1 U35 ( .A(a[12]), .B(n24), .Y(n4) );
  XOR2X1 U36 ( .A(a[8]), .B(a[7]), .Y(n24) );
  XOR2X1 U37 ( .A(a[3]), .B(a[8]), .Y(n2) );
  XOR2X1 U38 ( .A(a[9]), .B(a[8]), .Y(n22) );
  XOR2X1 U39 ( .A(a[6]), .B(a[1]), .Y(n19) );
  XOR2X1 U40 ( .A(a[11]), .B(n13), .Y(n21) );
  XOR2X1 U41 ( .A(a[0]), .B(n6), .Y(n31) );
  XOR2X1 U42 ( .A(n20), .B(n21), .Y(c[2]) );
  XOR2X1 U43 ( .A(a[1]), .B(n22), .Y(n20) );
endmodule


module multiply_3967 ( a, c );
  input [12:0] a;
  output [12:0] c;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;

  XOR2X1 U1 ( .A(n8), .B(n20), .Y(c[1]) );
  XOR2X1 U2 ( .A(n13), .B(n14), .Y(c[5]) );
  XOR2X1 U3 ( .A(n3), .B(n17), .Y(n13) );
  XOR2X1 U4 ( .A(n15), .B(n16), .Y(n14) );
  XOR2X1 U5 ( .A(n8), .B(n9), .Y(n7) );
  XOR2X1 U6 ( .A(n3), .B(n12), .Y(n11) );
  XNOR2X1 U7 ( .A(n18), .B(n19), .Y(c[4]) );
  XNOR2X1 U8 ( .A(n20), .B(n9), .Y(n19) );
  XOR2X1 U9 ( .A(n8), .B(n12), .Y(c[3]) );
  XOR2X1 U10 ( .A(n5), .B(n8), .Y(c[11]) );
  XOR2X1 U11 ( .A(n10), .B(n11), .Y(c[6]) );
  XOR2X1 U12 ( .A(a[11]), .B(n1), .Y(n10) );
  XOR2X1 U13 ( .A(n6), .B(n7), .Y(c[7]) );
  XOR2X1 U14 ( .A(a[4]), .B(a[2]), .Y(n6) );
  XOR2X1 U15 ( .A(n15), .B(n22), .Y(c[12]) );
  XOR2X1 U16 ( .A(a[7]), .B(a[0]), .Y(n22) );
  XOR2X1 U17 ( .A(a[10]), .B(a[9]), .Y(n15) );
  XOR2X1 U18 ( .A(a[12]), .B(a[8]), .Y(n8) );
  XOR2X1 U19 ( .A(a[5]), .B(a[11]), .Y(n9) );
  XOR2X1 U20 ( .A(a[0]), .B(a[11]), .Y(n16) );
  XOR2X1 U21 ( .A(a[1]), .B(a[4]), .Y(n12) );
  XOR2X1 U22 ( .A(a[12]), .B(a[3]), .Y(n3) );
  XOR2X1 U23 ( .A(a[6]), .B(a[9]), .Y(n5) );
  XOR2X1 U24 ( .A(a[10]), .B(a[7]), .Y(n1) );
  XOR2X1 U25 ( .A(a[2]), .B(n15), .Y(n20) );
  XOR2X1 U26 ( .A(a[1]), .B(a[8]), .Y(n18) );
  XOR2X1 U27 ( .A(a[6]), .B(a[2]), .Y(n17) );
  XOR2X1 U28 ( .A(n18), .B(n24), .Y(c[0]) );
  XOR2X1 U29 ( .A(a[10]), .B(n16), .Y(n24) );
  XOR2X1 U30 ( .A(n15), .B(n21), .Y(c[2]) );
  XOR2X1 U31 ( .A(a[3]), .B(a[11]), .Y(n21) );
  XOR2X1 U32 ( .A(n3), .B(n4), .Y(c[8]) );
  XOR2X1 U33 ( .A(a[5]), .B(n5), .Y(n4) );
  XOR2X1 U34 ( .A(n1), .B(n2), .Y(c[9]) );
  XOR2X1 U35 ( .A(a[6]), .B(a[4]), .Y(n2) );
  XOR2X1 U36 ( .A(n9), .B(n23), .Y(c[10]) );
  XOR2X1 U37 ( .A(a[8]), .B(a[7]), .Y(n23) );
endmodule


module mux_13_53 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n1, n2;

  BUFX3 U1 ( .A(n17), .Y(n2) );
  INVX1 U2 ( .A(n1), .Y(n17) );
  BUFX3 U3 ( .A(sel), .Y(n1) );
  INVX1 U4 ( .A(n29), .Y(out[0]) );
  AOI22X1 U5 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n2), .Y(n29) );
  INVX1 U6 ( .A(n25), .Y(out[1]) );
  AOI22X1 U7 ( .A0(a[1]), .A1(n1), .B0(b[1]), .B1(n17), .Y(n25) );
  INVX1 U8 ( .A(n24), .Y(out[2]) );
  AOI22X1 U9 ( .A0(a[2]), .A1(n1), .B0(b[2]), .B1(n2), .Y(n24) );
  INVX1 U10 ( .A(n23), .Y(out[3]) );
  AOI22X1 U11 ( .A0(a[3]), .A1(n1), .B0(b[3]), .B1(n2), .Y(n23) );
  INVX1 U12 ( .A(n22), .Y(out[4]) );
  AOI22X1 U13 ( .A0(a[4]), .A1(n1), .B0(b[4]), .B1(n2), .Y(n22) );
  INVX1 U14 ( .A(n21), .Y(out[5]) );
  AOI22X1 U15 ( .A0(a[5]), .A1(n1), .B0(b[5]), .B1(n2), .Y(n21) );
  INVX1 U16 ( .A(n20), .Y(out[6]) );
  AOI22X1 U17 ( .A0(a[6]), .A1(n1), .B0(b[6]), .B1(n2), .Y(n20) );
  INVX1 U18 ( .A(n19), .Y(out[7]) );
  AOI22X1 U19 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n2), .Y(n19) );
  INVX1 U20 ( .A(n18), .Y(out[8]) );
  AOI22X1 U21 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n2), .Y(n18) );
  INVX1 U22 ( .A(n16), .Y(out[9]) );
  AOI22X1 U23 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n16) );
  INVX1 U24 ( .A(n28), .Y(out[10]) );
  AOI22X1 U25 ( .A0(a[10]), .A1(sel), .B0(b[10]), .B1(n17), .Y(n28) );
  INVX1 U26 ( .A(n27), .Y(out[11]) );
  AOI22X1 U27 ( .A0(a[11]), .A1(n1), .B0(b[11]), .B1(n17), .Y(n27) );
  INVX1 U28 ( .A(n26), .Y(out[12]) );
  AOI22X1 U29 ( .A0(a[12]), .A1(sel), .B0(b[12]), .B1(n2), .Y(n26) );
endmodule


module feedback_ckt_16 ( Din, start, Qout, clk, reset );
  input [12:0] Din;
  output [12:0] Qout;
  input start, clk, reset;

  wire   [12:0] out;

  mux_13_20 mux ( .a(Qout), .b(Din), .sel(start), .out(out) );
  DFFRHQX1 \D_reg[0]  ( .D(out[0]), .CK(clk), .RN(reset), .Q(Qout[0]) );
  DFFRHQX1 \D_reg[1]  ( .D(out[1]), .CK(clk), .RN(reset), .Q(Qout[1]) );
  DFFRHQX1 \D_reg[4]  ( .D(out[4]), .CK(clk), .RN(reset), .Q(Qout[4]) );
  DFFRHQX1 \D_reg[10]  ( .D(out[10]), .CK(clk), .RN(reset), .Q(Qout[10]) );
  DFFRHQX1 \D_reg[2]  ( .D(out[2]), .CK(clk), .RN(reset), .Q(Qout[2]) );
  DFFRHQX1 \D_reg[5]  ( .D(out[5]), .CK(clk), .RN(reset), .Q(Qout[5]) );
  DFFRHQX1 \D_reg[11]  ( .D(out[11]), .CK(clk), .RN(reset), .Q(Qout[11]) );
  DFFRHQX1 \D_reg[3]  ( .D(out[3]), .CK(clk), .RN(reset), .Q(Qout[3]) );
  DFFRHQX1 \D_reg[12]  ( .D(out[12]), .CK(clk), .RN(reset), .Q(Qout[12]) );
  DFFRHQX1 \D_reg[9]  ( .D(out[9]), .CK(clk), .RN(reset), .Q(Qout[9]) );
  DFFRHQX1 \D_reg[7]  ( .D(out[7]), .CK(clk), .RN(reset), .Q(Qout[7]) );
  DFFRHQX1 \D_reg[8]  ( .D(out[8]), .CK(clk), .RN(reset), .Q(Qout[8]) );
  DFFRHQX1 \D_reg[6]  ( .D(out[6]), .CK(clk), .RN(reset), .Q(Qout[6]) );
endmodule


module euclidean_cell_3 ( deg_Ri, deg_Qi, stop_i, Rin, Qin, Lin, Uin, start, 
        start_cnt, deg_Ro, deg_Qo, stop_o, Rout, Qout, Lout, Uout, st_out, clk, 
        reset );
  input [4:0] deg_Ri;
  input [4:0] deg_Qi;
  input [12:0] Rin;
  input [12:0] Qin;
  input [12:0] Lin;
  input [12:0] Uin;
  output [4:0] deg_Ro;
  output [4:0] deg_Qo;
  output [12:0] Rout;
  output [12:0] Qout;
  output [12:0] Lout;
  output [12:0] Uout;
  input stop_i, start, start_cnt, clk, reset;
  output stop_o, st_out;
  wire   sw, start_temp, S2, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n135, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n2, n136, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309;
  wire   [12:0] d1out;
  wire   [12:0] Q1;
  wire   [12:0] R1;
  wire   [12:0] r_mux;
  wire   [12:0] q_mux;
  wire   [12:0] U1;
  wire   [12:0] L1;
  wire   [12:0] l_mux;
  wire   [12:0] u_mux;
  wire   [12:0] d2out;
  wire   [12:0] d3out;
  wire   [12:0] d4out;
  wire   [12:0] R2;
  wire   [12:0] m1out;
  wire   [12:0] Q2;
  wire   [12:0] m2out;
  wire   [12:0] L2;
  wire   [12:0] m3out;
  wire   [12:0] U2;
  wire   [12:0] m4out;
  wire   [12:0] add1out;
  wire   [12:0] add2out;
  wire   [12:0] Q3;
  wire   [12:0] U3;

  DFFRHQX4 \R2_reg[11]  ( .D(n217), .CK(clk), .RN(reset), .Q(R2[11]) );
  DFFRHQX4 \U2_reg[10]  ( .D(n166), .CK(clk), .RN(reset), .Q(U2[10]) );
  DFFRHQX4 \U2_reg[11]  ( .D(n165), .CK(clk), .RN(reset), .Q(U2[11]) );
  DFFRHQX4 \L2_reg[12]  ( .D(n151), .CK(clk), .RN(reset), .Q(L2[12]) );
  degree_computation_3 degree1 ( .deg_Ri(deg_Ri), .deg_Qi(deg_Qi), .stop_i(
        n270), .d1out(d1out), .start(start), .deg_Ro(deg_Ro), .deg_Qo(deg_Qo), 
        .stop_o(stop_o), .sw(sw), .clk(clk), .reset(reset) );
  mux_13_52 m1 ( .a(Q1), .b(R1), .sel(sw), .out(r_mux) );
  mux_13_51 m2 ( .a(R1), .b(Q1), .sel(sw), .out(q_mux) );
  mux_13_50 m3 ( .a(U1), .b(L1), .sel(sw), .out(l_mux) );
  mux_13_49 m4 ( .a(L1), .b(U1), .sel(sw), .out(u_mux) );
  feedback_ckt_15 D1 ( .Din(q_mux), .start(start_temp), .Qout(d1out), .clk(clk), .reset(reset) );
  feedback_ckt_14 D2 ( .Din(r_mux), .start(start_temp), .Qout(d2out), .clk(clk), .reset(reset) );
  feedback_ckt_13 D3 ( .Din(q_mux), .start(start_temp), .Qout(d3out), .clk(clk), .reset(reset) );
  feedback_ckt_12 D4 ( .Din(r_mux), .start(n136), .Qout(d4out), .clk(clk), 
        .reset(reset) );
  multiplier_15 mx1 ( .a(R2), .b(d1out), .c(m1out) );
  multiplier_14 mx2 ( .a(d2out), .b(Q2), .c(m2out) );
  multiplier_13 mx3 ( .a(L2), .b(d3out), .c(m3out) );
  multiplier_12 mx4 ( .a(d4out), .b(U2), .c(m4out) );
  mux_13_48 m5 ( .a(R2), .b(add1out), .sel(n270), .out(Rout) );
  mux_13_47 m6 ( .a(Q2), .b(Q3), .sel(n270), .out(Qout) );
  mux_13_46 m7 ( .a(L2), .b(add2out), .sel(n270), .out(Lout) );
  mux_13_45 m8 ( .a(U2), .b(U3), .sel(n270), .out(Uout) );
  DFFSX1 S3_reg ( .D(n137), .CK(clk), .SN(reset), .Q(st_out), .QN(n135) );
  DFFSX1 S2_reg ( .D(n268), .CK(clk), .SN(reset), .Q(S2) );
  DFFRHQX1 \Q3_reg[12]  ( .D(n215), .CK(clk), .RN(reset), .Q(Q3[12]) );
  DFFRHQX1 \Q3_reg[11]  ( .D(n214), .CK(clk), .RN(reset), .Q(Q3[11]) );
  DFFRHQX1 \Q3_reg[10]  ( .D(n213), .CK(clk), .RN(reset), .Q(Q3[10]) );
  DFFRHQX1 \Q3_reg[9]  ( .D(n212), .CK(clk), .RN(reset), .Q(Q3[9]) );
  DFFRHQX1 \Q3_reg[8]  ( .D(n211), .CK(clk), .RN(reset), .Q(Q3[8]) );
  DFFRHQX1 \Q3_reg[7]  ( .D(n210), .CK(clk), .RN(reset), .Q(Q3[7]) );
  DFFRHQX1 \Q3_reg[6]  ( .D(n209), .CK(clk), .RN(reset), .Q(Q3[6]) );
  DFFRHQX1 \Q3_reg[5]  ( .D(n208), .CK(clk), .RN(reset), .Q(Q3[5]) );
  DFFRHQX1 \Q3_reg[4]  ( .D(n207), .CK(clk), .RN(reset), .Q(Q3[4]) );
  DFFRHQX1 \Q3_reg[3]  ( .D(n206), .CK(clk), .RN(reset), .Q(Q3[3]) );
  DFFRHQX1 \Q3_reg[2]  ( .D(n205), .CK(clk), .RN(reset), .Q(Q3[2]) );
  DFFRHQX1 \Q3_reg[1]  ( .D(n204), .CK(clk), .RN(reset), .Q(Q3[1]) );
  DFFRHQX1 \Q3_reg[0]  ( .D(n203), .CK(clk), .RN(reset), .Q(Q3[0]) );
  DFFRHQX1 \U3_reg[12]  ( .D(n150), .CK(clk), .RN(reset), .Q(U3[12]) );
  DFFRHQX1 \U3_reg[11]  ( .D(n149), .CK(clk), .RN(reset), .Q(U3[11]) );
  DFFRHQX1 \U3_reg[10]  ( .D(n148), .CK(clk), .RN(reset), .Q(U3[10]) );
  DFFRHQX1 \U3_reg[9]  ( .D(n147), .CK(clk), .RN(reset), .Q(U3[9]) );
  DFFRHQX1 \U3_reg[8]  ( .D(n146), .CK(clk), .RN(reset), .Q(U3[8]) );
  DFFRHQX1 \U3_reg[7]  ( .D(n145), .CK(clk), .RN(reset), .Q(U3[7]) );
  DFFRHQX1 \U3_reg[6]  ( .D(n144), .CK(clk), .RN(reset), .Q(U3[6]) );
  DFFRHQX1 \U3_reg[5]  ( .D(n143), .CK(clk), .RN(reset), .Q(U3[5]) );
  DFFRHQX1 \U3_reg[4]  ( .D(n142), .CK(clk), .RN(reset), .Q(U3[4]) );
  DFFRHQX1 \U3_reg[3]  ( .D(n141), .CK(clk), .RN(reset), .Q(U3[3]) );
  DFFRHQX1 \U3_reg[2]  ( .D(n140), .CK(clk), .RN(reset), .Q(U3[2]) );
  DFFRHQX1 \U3_reg[1]  ( .D(n139), .CK(clk), .RN(reset), .Q(U3[1]) );
  DFFRHQX1 \U3_reg[0]  ( .D(n138), .CK(clk), .RN(reset), .Q(U3[0]) );
  DFFRHQX1 \R1_reg[12]  ( .D(n267), .CK(clk), .RN(reset), .Q(R1[12]) );
  DFFRHQX1 \R1_reg[11]  ( .D(n266), .CK(clk), .RN(reset), .Q(R1[11]) );
  DFFRHQX1 \R1_reg[10]  ( .D(n265), .CK(clk), .RN(reset), .Q(R1[10]) );
  DFFRHQX1 \R1_reg[8]  ( .D(n263), .CK(clk), .RN(reset), .Q(R1[8]) );
  DFFRHQX1 \R1_reg[7]  ( .D(n262), .CK(clk), .RN(reset), .Q(R1[7]) );
  DFFRHQX1 \R1_reg[6]  ( .D(n261), .CK(clk), .RN(reset), .Q(R1[6]) );
  DFFRHQX1 \R1_reg[5]  ( .D(n260), .CK(clk), .RN(reset), .Q(R1[5]) );
  DFFRHQX1 \R1_reg[4]  ( .D(n259), .CK(clk), .RN(reset), .Q(R1[4]) );
  DFFRHQX1 \R1_reg[3]  ( .D(n258), .CK(clk), .RN(reset), .Q(R1[3]) );
  DFFRHQX1 \R1_reg[2]  ( .D(n257), .CK(clk), .RN(reset), .Q(R1[2]) );
  DFFRHQX1 \R1_reg[1]  ( .D(n256), .CK(clk), .RN(reset), .Q(R1[1]) );
  DFFRHQX1 \R1_reg[0]  ( .D(n255), .CK(clk), .RN(reset), .Q(R1[0]) );
  DFFRHQX1 \Q1_reg[12]  ( .D(n254), .CK(clk), .RN(reset), .Q(Q1[12]) );
  DFFRHQX1 \Q1_reg[11]  ( .D(n253), .CK(clk), .RN(reset), .Q(Q1[11]) );
  DFFRHQX1 \Q1_reg[10]  ( .D(n252), .CK(clk), .RN(reset), .Q(Q1[10]) );
  DFFRHQX1 \Q1_reg[8]  ( .D(n250), .CK(clk), .RN(reset), .Q(Q1[8]) );
  DFFRHQX1 \Q1_reg[7]  ( .D(n249), .CK(clk), .RN(reset), .Q(Q1[7]) );
  DFFRHQX1 \Q1_reg[6]  ( .D(n248), .CK(clk), .RN(reset), .Q(Q1[6]) );
  DFFRHQX1 \Q1_reg[5]  ( .D(n247), .CK(clk), .RN(reset), .Q(Q1[5]) );
  DFFRHQX1 \Q1_reg[4]  ( .D(n246), .CK(clk), .RN(reset), .Q(Q1[4]) );
  DFFRHQX1 \Q1_reg[3]  ( .D(n245), .CK(clk), .RN(reset), .Q(Q1[3]) );
  DFFRHQX1 \Q1_reg[2]  ( .D(n244), .CK(clk), .RN(reset), .Q(Q1[2]) );
  DFFRHQX1 \Q1_reg[1]  ( .D(n243), .CK(clk), .RN(reset), .Q(Q1[1]) );
  DFFRHQX1 \Q1_reg[0]  ( .D(n242), .CK(clk), .RN(reset), .Q(Q1[0]) );
  DFFRHQX1 \L1_reg[12]  ( .D(n202), .CK(clk), .RN(reset), .Q(L1[12]) );
  DFFRHQX1 \L1_reg[11]  ( .D(n201), .CK(clk), .RN(reset), .Q(L1[11]) );
  DFFRHQX1 \L1_reg[10]  ( .D(n200), .CK(clk), .RN(reset), .Q(L1[10]) );
  DFFRHQX1 \L1_reg[8]  ( .D(n198), .CK(clk), .RN(reset), .Q(L1[8]) );
  DFFRHQX1 \L1_reg[7]  ( .D(n197), .CK(clk), .RN(reset), .Q(L1[7]) );
  DFFRHQX1 \L1_reg[6]  ( .D(n196), .CK(clk), .RN(reset), .Q(L1[6]) );
  DFFRHQX1 \L1_reg[5]  ( .D(n195), .CK(clk), .RN(reset), .Q(L1[5]) );
  DFFRHQX1 \L1_reg[4]  ( .D(n194), .CK(clk), .RN(reset), .Q(L1[4]) );
  DFFRHQX1 \L1_reg[3]  ( .D(n193), .CK(clk), .RN(reset), .Q(L1[3]) );
  DFFRHQX1 \L1_reg[2]  ( .D(n192), .CK(clk), .RN(reset), .Q(L1[2]) );
  DFFRHQX1 \L1_reg[1]  ( .D(n191), .CK(clk), .RN(reset), .Q(L1[1]) );
  DFFRHQX1 \L1_reg[0]  ( .D(n190), .CK(clk), .RN(reset), .Q(L1[0]) );
  DFFRHQX1 \U1_reg[12]  ( .D(n189), .CK(clk), .RN(reset), .Q(U1[12]) );
  DFFRHQX1 \U1_reg[11]  ( .D(n188), .CK(clk), .RN(reset), .Q(U1[11]) );
  DFFRHQX1 \U1_reg[10]  ( .D(n187), .CK(clk), .RN(reset), .Q(U1[10]) );
  DFFRHQX1 \U1_reg[8]  ( .D(n185), .CK(clk), .RN(reset), .Q(U1[8]) );
  DFFRHQX1 \U1_reg[7]  ( .D(n184), .CK(clk), .RN(reset), .Q(U1[7]) );
  DFFRHQX1 \U1_reg[6]  ( .D(n183), .CK(clk), .RN(reset), .Q(U1[6]) );
  DFFRHQX1 \U1_reg[5]  ( .D(n182), .CK(clk), .RN(reset), .Q(U1[5]) );
  DFFRHQX1 \U1_reg[4]  ( .D(n181), .CK(clk), .RN(reset), .Q(U1[4]) );
  DFFRHQX1 \U1_reg[3]  ( .D(n180), .CK(clk), .RN(reset), .Q(U1[3]) );
  DFFRHQX1 \U1_reg[2]  ( .D(n179), .CK(clk), .RN(reset), .Q(U1[2]) );
  DFFRHQX1 \U1_reg[1]  ( .D(n178), .CK(clk), .RN(reset), .Q(U1[1]) );
  DFFRHQX1 \U1_reg[0]  ( .D(n177), .CK(clk), .RN(reset), .Q(U1[0]) );
  DFFRHQX1 \R1_reg[9]  ( .D(n264), .CK(clk), .RN(reset), .Q(R1[9]) );
  DFFRHQX1 \Q1_reg[9]  ( .D(n251), .CK(clk), .RN(reset), .Q(Q1[9]) );
  DFFRHQX1 \L1_reg[9]  ( .D(n199), .CK(clk), .RN(reset), .Q(L1[9]) );
  DFFRHQX1 \U1_reg[9]  ( .D(n186), .CK(clk), .RN(reset), .Q(U1[9]) );
  DFFSX1 S1_reg ( .D(n269), .CK(clk), .SN(reset), .Q(start_temp), .QN(n2) );
  DFFRHQX1 \R2_reg[0]  ( .D(n228), .CK(clk), .RN(reset), .Q(R2[0]) );
  DFFRHQX1 \R2_reg[1]  ( .D(n227), .CK(clk), .RN(reset), .Q(R2[1]) );
  DFFRHQX1 \R2_reg[2]  ( .D(n226), .CK(clk), .RN(reset), .Q(R2[2]) );
  DFFRHQX1 \R2_reg[6]  ( .D(n222), .CK(clk), .RN(reset), .Q(R2[6]) );
  DFFRHQX1 \L2_reg[0]  ( .D(n163), .CK(clk), .RN(reset), .Q(L2[0]) );
  DFFRHQX1 \L2_reg[1]  ( .D(n162), .CK(clk), .RN(reset), .Q(L2[1]) );
  DFFRHQX1 \L2_reg[2]  ( .D(n161), .CK(clk), .RN(reset), .Q(L2[2]) );
  DFFRHQX1 \L2_reg[6]  ( .D(n157), .CK(clk), .RN(reset), .Q(L2[6]) );
  DFFRHQX1 \R2_reg[3]  ( .D(n225), .CK(clk), .RN(reset), .Q(R2[3]) );
  DFFRHQX1 \R2_reg[4]  ( .D(n224), .CK(clk), .RN(reset), .Q(R2[4]) );
  DFFRHQX1 \R2_reg[7]  ( .D(n221), .CK(clk), .RN(reset), .Q(R2[7]) );
  DFFRHQX1 \R2_reg[8]  ( .D(n220), .CK(clk), .RN(reset), .Q(R2[8]) );
  DFFRHQX1 \R2_reg[9]  ( .D(n219), .CK(clk), .RN(reset), .Q(R2[9]) );
  DFFRHQX1 \R2_reg[10]  ( .D(n218), .CK(clk), .RN(reset), .Q(R2[10]) );
  DFFRHQX1 \L2_reg[3]  ( .D(n160), .CK(clk), .RN(reset), .Q(L2[3]) );
  DFFRHQX1 \L2_reg[4]  ( .D(n159), .CK(clk), .RN(reset), .Q(L2[4]) );
  DFFRHQX1 \L2_reg[5]  ( .D(n158), .CK(clk), .RN(reset), .Q(L2[5]) );
  DFFRHQX1 \L2_reg[7]  ( .D(n156), .CK(clk), .RN(reset), .Q(L2[7]) );
  DFFRHQX1 \L2_reg[8]  ( .D(n155), .CK(clk), .RN(reset), .Q(L2[8]) );
  DFFRHQX1 \L2_reg[9]  ( .D(n154), .CK(clk), .RN(reset), .Q(L2[9]) );
  DFFRHQX1 \L2_reg[10]  ( .D(n153), .CK(clk), .RN(reset), .Q(L2[10]) );
  DFFRHQX1 \Q2_reg[2]  ( .D(n239), .CK(clk), .RN(reset), .Q(Q2[2]) );
  DFFRHQX1 \Q2_reg[6]  ( .D(n235), .CK(clk), .RN(reset), .Q(Q2[6]) );
  DFFRHQX1 \Q2_reg[7]  ( .D(n234), .CK(clk), .RN(reset), .Q(Q2[7]) );
  DFFRHQX1 \Q2_reg[12]  ( .D(n229), .CK(clk), .RN(reset), .Q(Q2[12]) );
  DFFRHQX1 \U2_reg[2]  ( .D(n174), .CK(clk), .RN(reset), .Q(U2[2]) );
  DFFRHQX1 \U2_reg[5]  ( .D(n171), .CK(clk), .RN(reset), .Q(U2[5]) );
  DFFRHQX1 \U2_reg[6]  ( .D(n170), .CK(clk), .RN(reset), .Q(U2[6]) );
  DFFRHQX1 \U2_reg[7]  ( .D(n169), .CK(clk), .RN(reset), .Q(U2[7]) );
  DFFRHQX1 \U2_reg[8]  ( .D(n168), .CK(clk), .RN(reset), .Q(U2[8]) );
  DFFRHQX1 \U2_reg[12]  ( .D(n164), .CK(clk), .RN(reset), .Q(U2[12]) );
  DFFRHQX1 \U2_reg[9]  ( .D(n167), .CK(clk), .RN(reset), .Q(U2[9]) );
  DFFRHQX1 \Q2_reg[0]  ( .D(n241), .CK(clk), .RN(reset), .Q(Q2[0]) );
  DFFRHQX1 \U2_reg[0]  ( .D(n176), .CK(clk), .RN(reset), .Q(U2[0]) );
  DFFRHQX1 \Q2_reg[1]  ( .D(n240), .CK(clk), .RN(reset), .Q(Q2[1]) );
  DFFRHQX1 \U2_reg[1]  ( .D(n175), .CK(clk), .RN(reset), .Q(U2[1]) );
  DFFRHQX2 \Q2_reg[4]  ( .D(n237), .CK(clk), .RN(reset), .Q(Q2[4]) );
  DFFRHQX2 \U2_reg[4]  ( .D(n172), .CK(clk), .RN(reset), .Q(U2[4]) );
  DFFRHQX2 \L2_reg[11]  ( .D(n152), .CK(clk), .RN(reset), .Q(L2[11]) );
  DFFRHQX2 \Q2_reg[5]  ( .D(n236), .CK(clk), .RN(reset), .Q(Q2[5]) );
  DFFRHQX1 \Q2_reg[8]  ( .D(n233), .CK(clk), .RN(reset), .Q(Q2[8]) );
  DFFRHQX1 \Q2_reg[9]  ( .D(n232), .CK(clk), .RN(reset), .Q(Q2[9]) );
  DFFRHQX2 \U2_reg[3]  ( .D(n173), .CK(clk), .RN(reset), .Q(U2[3]) );
  DFFRHQX2 \Q2_reg[3]  ( .D(n238), .CK(clk), .RN(reset), .Q(Q2[3]) );
  DFFRHQX2 \Q2_reg[10]  ( .D(n231), .CK(clk), .RN(reset), .Q(Q2[10]) );
  DFFRHQX2 \R2_reg[12]  ( .D(n216), .CK(clk), .RN(reset), .Q(R2[12]) );
  DFFRHQX1 \R2_reg[5]  ( .D(n223), .CK(clk), .RN(reset), .Q(R2[5]) );
  DFFRHQX4 \Q2_reg[11]  ( .D(n230), .CK(clk), .RN(reset), .Q(Q2[11]) );
  AOI22XL U2_inst ( .A0(n291), .A1(U2[2]), .B0(u_mux[2]), .B1(n283), .Y(n38)
         );
  AOI22XL U3_inst ( .A0(n273), .A1(U2[2]), .B0(U3[2]), .B1(n304), .Y(n4) );
  XOR2X1 U4 ( .A(m2out[4]), .B(m1out[4]), .Y(add1out[4]) );
  XOR2X1 U5 ( .A(m4out[4]), .B(m3out[4]), .Y(add2out[4]) );
  XOR2X1 U6 ( .A(m4out[8]), .B(m3out[8]), .Y(add2out[8]) );
  XOR2X1 U7 ( .A(m4out[11]), .B(m3out[11]), .Y(add2out[11]) );
  XOR2X1 U8 ( .A(m2out[5]), .B(m1out[5]), .Y(add1out[5]) );
  XOR2X1 U9 ( .A(m4out[5]), .B(m3out[5]), .Y(add2out[5]) );
  AOI22XL U10 ( .A0(R2[11]), .A1(n309), .B0(r_mux[11]), .B1(n286), .Y(n81) );
  AOI22XL U11 ( .A0(n278), .A1(U2[1]), .B0(U3[1]), .B1(n297), .Y(n3) );
  AOI22XL U12 ( .A0(n273), .A1(U2[3]), .B0(U3[3]), .B1(n294), .Y(n5) );
  AOI22XL U13 ( .A0(n276), .A1(U2[4]), .B0(U3[4]), .B1(n303), .Y(n6) );
  AOI22XL U14 ( .A0(n278), .A1(U2[5]), .B0(U3[5]), .B1(n293), .Y(n7) );
  AOI22XL U15 ( .A0(n274), .A1(U2[6]), .B0(U3[6]), .B1(n303), .Y(n8) );
  AOI22XL U16 ( .A0(n275), .A1(U2[7]), .B0(U3[7]), .B1(n295), .Y(n9) );
  AOI22XL U17 ( .A0(n275), .A1(U2[8]), .B0(U3[8]), .B1(n291), .Y(n10) );
  AOI22XL U18 ( .A0(n273), .A1(U2[9]), .B0(U3[9]), .B1(n295), .Y(n11) );
  AOI22XL U19 ( .A0(n276), .A1(U2[10]), .B0(U3[10]), .B1(n297), .Y(n12) );
  AOI22XL U20 ( .A0(n278), .A1(U2[11]), .B0(U3[11]), .B1(n293), .Y(n13) );
  AOI22XL U21 ( .A0(n276), .A1(U2[12]), .B0(U3[12]), .B1(n294), .Y(n14) );
  AOI22XL U22 ( .A0(n276), .A1(Q2[0]), .B0(Q3[0]), .B1(n296), .Y(n67) );
  AOI22XL U23 ( .A0(n277), .A1(Q2[1]), .B0(Q3[1]), .B1(n297), .Y(n68) );
  AOI22XL U24 ( .A0(n277), .A1(Q2[3]), .B0(Q3[3]), .B1(n297), .Y(n70) );
  AOI22XL U25 ( .A0(n278), .A1(Q2[5]), .B0(Q3[5]), .B1(n298), .Y(n72) );
  AOI22XL U26 ( .A0(n274), .A1(Q2[6]), .B0(Q3[6]), .B1(n293), .Y(n73) );
  AOI22XL U27 ( .A0(n277), .A1(Q2[9]), .B0(Q3[9]), .B1(n294), .Y(n76) );
  AOI22XL U28 ( .A0(n277), .A1(Q2[12]), .B0(Q3[12]), .B1(n296), .Y(n79) );
  AOI22XL U29 ( .A0(n308), .A1(U2[1]), .B0(u_mux[1]), .B1(n283), .Y(n39) );
  AOI22XL U30 ( .A0(n299), .A1(Q2[1]), .B0(q_mux[1]), .B1(n283), .Y(n104) );
  AOI22XL U31 ( .A0(n308), .A1(U2[11]), .B0(u_mux[11]), .B1(n286), .Y(n29) );
  AOI22XL U32 ( .A0(n298), .A1(U2[10]), .B0(u_mux[10]), .B1(n286), .Y(n30) );
  AOI22XL U33 ( .A0(n309), .A1(U2[3]), .B0(u_mux[3]), .B1(n306), .Y(n37) );
  AOI22XL U34 ( .A0(n293), .A1(Q2[11]), .B0(q_mux[11]), .B1(n306), .Y(n94) );
  AOI22XL U35 ( .A0(n308), .A1(Q2[10]), .B0(q_mux[10]), .B1(n288), .Y(n95) );
  AOI22XL U36 ( .A0(n296), .A1(Q2[3]), .B0(q_mux[3]), .B1(n287), .Y(n102) );
  AOI22XL U37 ( .A0(L2[12]), .A1(n294), .B0(l_mux[12]), .B1(n288), .Y(n15) );
  AOI22XL U38 ( .A0(R2[12]), .A1(n309), .B0(r_mux[12]), .B1(n285), .Y(n80) );
  AOI22XL U39 ( .A0(n274), .A1(Q2[4]), .B0(Q3[4]), .B1(n295), .Y(n71) );
  AOI22XL U40 ( .A0(n278), .A1(Q2[7]), .B0(Q3[7]), .B1(n309), .Y(n74) );
  AOI22XL U41 ( .A0(n274), .A1(Q2[8]), .B0(Q3[8]), .B1(n298), .Y(n75) );
  AOI22XL U42 ( .A0(n275), .A1(Q2[10]), .B0(Q3[10]), .B1(n295), .Y(n77) );
  AOI22XL U43 ( .A0(n277), .A1(Q2[11]), .B0(Q3[11]), .B1(n295), .Y(n78) );
  AOI22XL U44 ( .A0(n304), .A1(Q2[0]), .B0(q_mux[0]), .B1(n287), .Y(n105) );
  AOI22XL U45 ( .A0(n303), .A1(U2[8]), .B0(u_mux[8]), .B1(n284), .Y(n32) );
  AOI22XL U46 ( .A0(n292), .A1(U2[5]), .B0(u_mux[5]), .B1(n284), .Y(n35) );
  AOI22XL U47 ( .A0(n295), .A1(U2[0]), .B0(u_mux[0]), .B1(n287), .Y(n40) );
  AOI22XL U48 ( .A0(n291), .A1(Q2[12]), .B0(q_mux[12]), .B1(n285), .Y(n93) );
  AOI22XL U49 ( .A0(n303), .A1(Q2[9]), .B0(q_mux[9]), .B1(n283), .Y(n96) );
  AOI22XL U50 ( .A0(n295), .A1(Q2[8]), .B0(q_mux[8]), .B1(n284), .Y(n97) );
  AOI22XL U51 ( .A0(n303), .A1(Q2[7]), .B0(q_mux[7]), .B1(n285), .Y(n98) );
  AOI22XL U52 ( .A0(n294), .A1(Q2[6]), .B0(q_mux[6]), .B1(n305), .Y(n99) );
  AOI22XL U53 ( .A0(n297), .A1(Q2[5]), .B0(q_mux[5]), .B1(n283), .Y(n100) );
  AOI22XL U54 ( .A0(n301), .A1(Q2[4]), .B0(q_mux[4]), .B1(n306), .Y(n101) );
  AOI22XL U55 ( .A0(n299), .A1(U2[12]), .B0(u_mux[12]), .B1(n287), .Y(n28) );
  AOI22XL U56 ( .A0(n302), .A1(U2[9]), .B0(u_mux[9]), .B1(n288), .Y(n31) );
  AOI22XL U57 ( .A0(n301), .A1(U2[7]), .B0(u_mux[7]), .B1(start_cnt), .Y(n33)
         );
  AOI22XL U58 ( .A0(n296), .A1(U2[6]), .B0(u_mux[6]), .B1(n285), .Y(n34) );
  AOI22XL U59 ( .A0(n300), .A1(U2[4]), .B0(u_mux[4]), .B1(n305), .Y(n36) );
  AOI22XL U60 ( .A0(L2[10]), .A1(n293), .B0(l_mux[10]), .B1(n306), .Y(n17) );
  AOI22XL U61 ( .A0(L2[9]), .A1(n299), .B0(l_mux[9]), .B1(n282), .Y(n18) );
  AOI22XL U62 ( .A0(L2[8]), .A1(n300), .B0(l_mux[8]), .B1(n287), .Y(n19) );
  AOI22XL U63 ( .A0(L2[5]), .A1(n301), .B0(l_mux[5]), .B1(n287), .Y(n22) );
  AOI22XL U64 ( .A0(L2[3]), .A1(n298), .B0(l_mux[3]), .B1(n288), .Y(n24) );
  AOI22XL U65 ( .A0(R2[9]), .A1(n291), .B0(r_mux[9]), .B1(n285), .Y(n83) );
  AOI22XL U66 ( .A0(R2[8]), .A1(n308), .B0(r_mux[8]), .B1(n282), .Y(n84) );
  AOI22XL U67 ( .A0(R2[6]), .A1(n292), .B0(r_mux[6]), .B1(n285), .Y(n86) );
  AOI22XL U68 ( .A0(R2[10]), .A1(n297), .B0(r_mux[10]), .B1(n284), .Y(n82) );
  AOI22XL U69 ( .A0(R2[7]), .A1(n291), .B0(r_mux[7]), .B1(n287), .Y(n85) );
  AOI22XL U70 ( .A0(R2[5]), .A1(n296), .B0(r_mux[5]), .B1(n285), .Y(n87) );
  AOI22XL U71 ( .A0(R2[4]), .A1(n302), .B0(r_mux[4]), .B1(n284), .Y(n88) );
  AOI22XL U72 ( .A0(R2[3]), .A1(n292), .B0(r_mux[3]), .B1(n284), .Y(n89) );
  AOI22XL U73 ( .A0(n284), .A1(U2[0]), .B0(U3[0]), .B1(n298), .Y(n1) );
  INVX1 U74 ( .A(n304), .Y(n272) );
  INVX1 U75 ( .A(n304), .Y(n273) );
  INVX1 U76 ( .A(n301), .Y(n276) );
  INVX1 U77 ( .A(n301), .Y(n275) );
  INVX1 U78 ( .A(n301), .Y(n274) );
  INVX1 U79 ( .A(n300), .Y(n278) );
  INVX1 U80 ( .A(n300), .Y(n277) );
  INVX1 U81 ( .A(n293), .Y(n290) );
  INVX1 U82 ( .A(n293), .Y(n289) );
  INVX1 U83 ( .A(n298), .Y(n285) );
  INVX1 U84 ( .A(n296), .Y(n284) );
  INVX1 U85 ( .A(n294), .Y(n286) );
  INVX1 U86 ( .A(n294), .Y(n287) );
  INVX1 U87 ( .A(n296), .Y(n283) );
  INVX1 U88 ( .A(n299), .Y(n281) );
  INVX1 U89 ( .A(n298), .Y(n282) );
  INVX1 U90 ( .A(n299), .Y(n280) );
  INVX1 U91 ( .A(n299), .Y(n279) );
  INVX1 U92 ( .A(n294), .Y(n288) );
  INVX1 U93 ( .A(n305), .Y(n291) );
  INVX1 U94 ( .A(n305), .Y(n292) );
  INVX1 U95 ( .A(n307), .Y(n293) );
  INVX1 U96 ( .A(n306), .Y(n301) );
  INVX1 U97 ( .A(n305), .Y(n302) );
  INVX1 U98 ( .A(n306), .Y(n300) );
  INVX1 U99 ( .A(n305), .Y(n303) );
  INVX1 U100 ( .A(n306), .Y(n295) );
  INVX1 U101 ( .A(n307), .Y(n297) );
  INVX1 U102 ( .A(n307), .Y(n296) );
  INVX1 U103 ( .A(n306), .Y(n299) );
  INVX1 U104 ( .A(n307), .Y(n298) );
  INVX1 U105 ( .A(n307), .Y(n294) );
  INVX1 U106 ( .A(n305), .Y(n304) );
  INVX1 U107 ( .A(n309), .Y(n305) );
  INVX1 U108 ( .A(n309), .Y(n306) );
  INVX1 U109 ( .A(n308), .Y(n307) );
  INVX1 U110 ( .A(start_cnt), .Y(n308) );
  INVX1 U111 ( .A(start_cnt), .Y(n309) );
  XOR2X1 U112 ( .A(m3out[10]), .B(m4out[10]), .Y(add2out[10]) );
  XOR2X1 U113 ( .A(m1out[10]), .B(m2out[10]), .Y(add1out[10]) );
  XOR2X1 U114 ( .A(m1out[8]), .B(m2out[8]), .Y(add1out[8]) );
  XOR2X1 U115 ( .A(m4out[6]), .B(m3out[6]), .Y(add2out[6]) );
  XOR2X1 U116 ( .A(m2out[6]), .B(m1out[6]), .Y(add1out[6]) );
  XOR2X1 U117 ( .A(m4out[2]), .B(m3out[2]), .Y(add2out[2]) );
  XOR2X1 U118 ( .A(m4out[1]), .B(m3out[1]), .Y(add2out[1]) );
  XOR2X1 U119 ( .A(m2out[1]), .B(m1out[1]), .Y(add1out[1]) );
  XOR2X1 U120 ( .A(m2out[2]), .B(m1out[2]), .Y(add1out[2]) );
  XOR2X1 U121 ( .A(m4out[12]), .B(m3out[12]), .Y(add2out[12]) );
  XOR2X1 U122 ( .A(m2out[12]), .B(m1out[12]), .Y(add1out[12]) );
  INVX1 U123 ( .A(n271), .Y(n270) );
  XOR2X1 U124 ( .A(m1out[7]), .B(m2out[7]), .Y(add1out[7]) );
  XOR2X1 U125 ( .A(m3out[7]), .B(m4out[7]), .Y(add2out[7]) );
  XOR2X1 U126 ( .A(m3out[3]), .B(m4out[3]), .Y(add2out[3]) );
  XOR2X1 U127 ( .A(m3out[9]), .B(m4out[9]), .Y(add2out[9]) );
  XOR2X1 U128 ( .A(m1out[3]), .B(m2out[3]), .Y(add1out[3]) );
  XOR2X1 U129 ( .A(m1out[9]), .B(m2out[9]), .Y(add1out[9]) );
  XOR2X1 U130 ( .A(m1out[11]), .B(m2out[11]), .Y(add1out[11]) );
  XOR2X1 U131 ( .A(m4out[0]), .B(m3out[0]), .Y(add2out[0]) );
  XOR2X1 U132 ( .A(m2out[0]), .B(m1out[0]), .Y(add1out[0]) );
  INVX1 U133 ( .A(stop_i), .Y(n271) );
  INVX1 U134 ( .A(n133), .Y(n269) );
  AOI22X1 U135 ( .A0(n297), .A1(n136), .B0(start), .B1(n288), .Y(n133) );
  INVX1 U136 ( .A(n2), .Y(n136) );
  INVX1 U137 ( .A(n17), .Y(n153) );
  OAI2BB2X1 U138 ( .B0(n272), .B1(n135), .A0N(S2), .A1N(n272), .Y(n137) );
  INVX1 U139 ( .A(n16), .Y(n152) );
  INVX1 U140 ( .A(n3), .Y(n139) );
  INVX1 U141 ( .A(n39), .Y(n175) );
  INVX1 U142 ( .A(n68), .Y(n204) );
  INVX1 U143 ( .A(n104), .Y(n240) );
  INVX1 U144 ( .A(n1), .Y(n138) );
  INVX1 U145 ( .A(n40), .Y(n176) );
  INVX1 U146 ( .A(n67), .Y(n203) );
  INVX1 U147 ( .A(n105), .Y(n241) );
  INVX1 U148 ( .A(n11), .Y(n147) );
  INVX1 U149 ( .A(n31), .Y(n167) );
  INVX1 U150 ( .A(n76), .Y(n212) );
  INVX1 U151 ( .A(n96), .Y(n232) );
  INVX1 U152 ( .A(n4), .Y(n140) );
  INVX1 U153 ( .A(n5), .Y(n141) );
  INVX1 U154 ( .A(n6), .Y(n142) );
  INVX1 U155 ( .A(n7), .Y(n143) );
  INVX1 U156 ( .A(n8), .Y(n144) );
  INVX1 U157 ( .A(n9), .Y(n145) );
  INVX1 U158 ( .A(n10), .Y(n146) );
  INVX1 U159 ( .A(n12), .Y(n148) );
  INVX1 U160 ( .A(n13), .Y(n149) );
  INVX1 U161 ( .A(n14), .Y(n150) );
  INVX1 U162 ( .A(n28), .Y(n164) );
  INVX1 U163 ( .A(n29), .Y(n165) );
  INVX1 U164 ( .A(n30), .Y(n166) );
  INVX1 U165 ( .A(n32), .Y(n168) );
  INVX1 U166 ( .A(n33), .Y(n169) );
  INVX1 U167 ( .A(n34), .Y(n170) );
  INVX1 U168 ( .A(n35), .Y(n171) );
  INVX1 U169 ( .A(n36), .Y(n172) );
  INVX1 U170 ( .A(n37), .Y(n173) );
  INVX1 U171 ( .A(n38), .Y(n174) );
  INVX1 U172 ( .A(n69), .Y(n205) );
  AOI22X1 U173 ( .A0(n275), .A1(Q2[2]), .B0(Q3[2]), .B1(n291), .Y(n69) );
  INVX1 U174 ( .A(n70), .Y(n206) );
  INVX1 U175 ( .A(n71), .Y(n207) );
  INVX1 U176 ( .A(n72), .Y(n208) );
  INVX1 U177 ( .A(n73), .Y(n209) );
  INVX1 U178 ( .A(n74), .Y(n210) );
  INVX1 U179 ( .A(n75), .Y(n211) );
  INVX1 U180 ( .A(n77), .Y(n213) );
  INVX1 U181 ( .A(n78), .Y(n214) );
  INVX1 U182 ( .A(n79), .Y(n215) );
  INVX1 U183 ( .A(n93), .Y(n229) );
  INVX1 U184 ( .A(n94), .Y(n230) );
  INVX1 U185 ( .A(n95), .Y(n231) );
  INVX1 U186 ( .A(n97), .Y(n233) );
  INVX1 U187 ( .A(n98), .Y(n234) );
  INVX1 U188 ( .A(n99), .Y(n235) );
  INVX1 U189 ( .A(n100), .Y(n236) );
  INVX1 U190 ( .A(n101), .Y(n237) );
  INVX1 U191 ( .A(n102), .Y(n238) );
  INVX1 U192 ( .A(n103), .Y(n239) );
  AOI22X1 U193 ( .A0(n302), .A1(Q2[2]), .B0(q_mux[2]), .B1(n282), .Y(n103) );
  INVX1 U194 ( .A(n15), .Y(n151) );
  INVX1 U195 ( .A(n18), .Y(n154) );
  INVX1 U196 ( .A(n19), .Y(n155) );
  INVX1 U197 ( .A(n20), .Y(n156) );
  AOI22X1 U198 ( .A0(L2[7]), .A1(n303), .B0(l_mux[7]), .B1(n286), .Y(n20) );
  INVX1 U199 ( .A(n21), .Y(n157) );
  AOI22X1 U200 ( .A0(L2[6]), .A1(n296), .B0(l_mux[6]), .B1(n289), .Y(n21) );
  INVX1 U201 ( .A(n22), .Y(n158) );
  INVX1 U202 ( .A(n23), .Y(n159) );
  AOI22X1 U203 ( .A0(L2[4]), .A1(n303), .B0(l_mux[4]), .B1(n290), .Y(n23) );
  INVX1 U204 ( .A(n24), .Y(n160) );
  INVX1 U205 ( .A(n25), .Y(n161) );
  AOI22X1 U206 ( .A0(L2[2]), .A1(n297), .B0(l_mux[2]), .B1(n286), .Y(n25) );
  INVX1 U207 ( .A(n26), .Y(n162) );
  AOI22X1 U208 ( .A0(L2[1]), .A1(n292), .B0(l_mux[1]), .B1(n283), .Y(n26) );
  INVX1 U209 ( .A(n27), .Y(n163) );
  AOI22X1 U210 ( .A0(L2[0]), .A1(n304), .B0(l_mux[0]), .B1(n283), .Y(n27) );
  INVX1 U211 ( .A(n41), .Y(n177) );
  AOI22X1 U212 ( .A0(U1[0]), .A1(n298), .B0(Uin[0]), .B1(n288), .Y(n41) );
  INVX1 U213 ( .A(n42), .Y(n178) );
  AOI22X1 U214 ( .A0(U1[1]), .A1(n303), .B0(Uin[1]), .B1(n289), .Y(n42) );
  INVX1 U215 ( .A(n43), .Y(n179) );
  AOI22X1 U216 ( .A0(U1[2]), .A1(n300), .B0(Uin[2]), .B1(n290), .Y(n43) );
  INVX1 U217 ( .A(n44), .Y(n180) );
  AOI22X1 U218 ( .A0(U1[3]), .A1(n308), .B0(Uin[3]), .B1(n288), .Y(n44) );
  INVX1 U219 ( .A(n45), .Y(n181) );
  AOI22X1 U220 ( .A0(U1[4]), .A1(n302), .B0(Uin[4]), .B1(n285), .Y(n45) );
  INVX1 U221 ( .A(n46), .Y(n182) );
  AOI22X1 U222 ( .A0(U1[5]), .A1(n295), .B0(Uin[5]), .B1(n289), .Y(n46) );
  INVX1 U223 ( .A(n47), .Y(n183) );
  AOI22X1 U224 ( .A0(U1[6]), .A1(n292), .B0(Uin[6]), .B1(n286), .Y(n47) );
  INVX1 U225 ( .A(n48), .Y(n184) );
  AOI22X1 U226 ( .A0(U1[7]), .A1(n309), .B0(Uin[7]), .B1(n287), .Y(n48) );
  INVX1 U227 ( .A(n49), .Y(n185) );
  AOI22X1 U228 ( .A0(U1[8]), .A1(n299), .B0(Uin[8]), .B1(n282), .Y(n49) );
  INVX1 U229 ( .A(n50), .Y(n186) );
  AOI22X1 U230 ( .A0(U1[9]), .A1(n309), .B0(Uin[9]), .B1(n284), .Y(n50) );
  INVX1 U231 ( .A(n51), .Y(n187) );
  AOI22X1 U232 ( .A0(U1[10]), .A1(n291), .B0(Uin[10]), .B1(n289), .Y(n51) );
  INVX1 U233 ( .A(n52), .Y(n188) );
  AOI22X1 U234 ( .A0(U1[11]), .A1(n300), .B0(Uin[11]), .B1(n306), .Y(n52) );
  INVX1 U235 ( .A(n53), .Y(n189) );
  AOI22X1 U236 ( .A0(U1[12]), .A1(n299), .B0(Uin[12]), .B1(n290), .Y(n53) );
  INVX1 U237 ( .A(n54), .Y(n190) );
  AOI22X1 U238 ( .A0(L1[0]), .A1(n302), .B0(Lin[0]), .B1(n282), .Y(n54) );
  INVX1 U239 ( .A(n55), .Y(n191) );
  AOI22X1 U240 ( .A0(L1[1]), .A1(n304), .B0(Lin[1]), .B1(n283), .Y(n55) );
  INVX1 U241 ( .A(n56), .Y(n192) );
  AOI22X1 U242 ( .A0(L1[2]), .A1(n303), .B0(Lin[2]), .B1(n305), .Y(n56) );
  INVX1 U243 ( .A(n57), .Y(n193) );
  AOI22X1 U244 ( .A0(L1[3]), .A1(n301), .B0(Lin[3]), .B1(n305), .Y(n57) );
  INVX1 U245 ( .A(n58), .Y(n194) );
  AOI22X1 U246 ( .A0(L1[4]), .A1(n292), .B0(Lin[4]), .B1(n287), .Y(n58) );
  INVX1 U247 ( .A(n59), .Y(n195) );
  AOI22X1 U248 ( .A0(L1[5]), .A1(n302), .B0(Lin[5]), .B1(n284), .Y(n59) );
  INVX1 U249 ( .A(n60), .Y(n196) );
  AOI22X1 U250 ( .A0(L1[6]), .A1(n304), .B0(Lin[6]), .B1(n289), .Y(n60) );
  INVX1 U251 ( .A(n61), .Y(n197) );
  AOI22X1 U252 ( .A0(L1[7]), .A1(n292), .B0(Lin[7]), .B1(n290), .Y(n61) );
  INVX1 U253 ( .A(n62), .Y(n198) );
  AOI22X1 U254 ( .A0(L1[8]), .A1(n309), .B0(Lin[8]), .B1(n290), .Y(n62) );
  INVX1 U255 ( .A(n63), .Y(n199) );
  AOI22X1 U256 ( .A0(L1[9]), .A1(n294), .B0(Lin[9]), .B1(n290), .Y(n63) );
  INVX1 U257 ( .A(n64), .Y(n200) );
  AOI22X1 U258 ( .A0(L1[10]), .A1(n293), .B0(Lin[10]), .B1(n289), .Y(n64) );
  INVX1 U259 ( .A(n65), .Y(n201) );
  AOI22X1 U260 ( .A0(L1[11]), .A1(n308), .B0(Lin[11]), .B1(n289), .Y(n65) );
  INVX1 U261 ( .A(n66), .Y(n202) );
  AOI22X1 U262 ( .A0(L1[12]), .A1(n302), .B0(Lin[12]), .B1(n288), .Y(n66) );
  INVX1 U263 ( .A(n80), .Y(n216) );
  INVX1 U264 ( .A(n81), .Y(n217) );
  INVX1 U265 ( .A(n82), .Y(n218) );
  INVX1 U266 ( .A(n83), .Y(n219) );
  INVX1 U267 ( .A(n84), .Y(n220) );
  INVX1 U268 ( .A(n85), .Y(n221) );
  INVX1 U269 ( .A(n86), .Y(n222) );
  INVX1 U270 ( .A(n87), .Y(n223) );
  INVX1 U271 ( .A(n88), .Y(n224) );
  INVX1 U272 ( .A(n89), .Y(n225) );
  INVX1 U273 ( .A(n90), .Y(n226) );
  AOI22X1 U274 ( .A0(R2[2]), .A1(n299), .B0(r_mux[2]), .B1(n290), .Y(n90) );
  INVX1 U275 ( .A(n91), .Y(n227) );
  AOI22X1 U276 ( .A0(R2[1]), .A1(n291), .B0(r_mux[1]), .B1(n286), .Y(n91) );
  INVX1 U277 ( .A(n92), .Y(n228) );
  AOI22X1 U278 ( .A0(R2[0]), .A1(n299), .B0(r_mux[0]), .B1(n289), .Y(n92) );
  INVX1 U279 ( .A(n106), .Y(n242) );
  AOI22X1 U280 ( .A0(Q1[0]), .A1(n304), .B0(Qin[0]), .B1(n284), .Y(n106) );
  INVX1 U281 ( .A(n107), .Y(n243) );
  AOI22X1 U282 ( .A0(Q1[1]), .A1(n302), .B0(Qin[1]), .B1(n282), .Y(n107) );
  INVX1 U283 ( .A(n108), .Y(n244) );
  AOI22X1 U284 ( .A0(Q1[2]), .A1(n301), .B0(Qin[2]), .B1(n287), .Y(n108) );
  INVX1 U285 ( .A(n109), .Y(n245) );
  AOI22X1 U286 ( .A0(Q1[3]), .A1(n303), .B0(Qin[3]), .B1(n288), .Y(n109) );
  INVX1 U287 ( .A(n110), .Y(n246) );
  AOI22X1 U288 ( .A0(Q1[4]), .A1(n291), .B0(Qin[4]), .B1(n289), .Y(n110) );
  INVX1 U289 ( .A(n111), .Y(n247) );
  AOI22X1 U290 ( .A0(Q1[5]), .A1(n300), .B0(Qin[5]), .B1(n283), .Y(n111) );
  INVX1 U291 ( .A(n112), .Y(n248) );
  AOI22X1 U292 ( .A0(Q1[6]), .A1(n301), .B0(Qin[6]), .B1(n286), .Y(n112) );
  INVX1 U293 ( .A(n113), .Y(n249) );
  AOI22X1 U294 ( .A0(Q1[7]), .A1(n300), .B0(Qin[7]), .B1(n286), .Y(n113) );
  INVX1 U295 ( .A(n114), .Y(n250) );
  AOI22X1 U296 ( .A0(Q1[8]), .A1(n297), .B0(Qin[8]), .B1(n290), .Y(n114) );
  INVX1 U297 ( .A(n115), .Y(n251) );
  AOI22X1 U298 ( .A0(Q1[9]), .A1(n304), .B0(Qin[9]), .B1(n282), .Y(n115) );
  INVX1 U299 ( .A(n116), .Y(n252) );
  AOI22X1 U300 ( .A0(Q1[10]), .A1(n309), .B0(Qin[10]), .B1(n282), .Y(n116) );
  INVX1 U301 ( .A(n117), .Y(n253) );
  AOI22X1 U302 ( .A0(Q1[11]), .A1(n302), .B0(Qin[11]), .B1(n290), .Y(n117) );
  INVX1 U303 ( .A(n118), .Y(n254) );
  AOI22X1 U304 ( .A0(Q1[12]), .A1(n296), .B0(Qin[12]), .B1(n281), .Y(n118) );
  INVX1 U305 ( .A(n119), .Y(n255) );
  AOI22X1 U306 ( .A0(R1[0]), .A1(n294), .B0(Rin[0]), .B1(n305), .Y(n119) );
  INVX1 U307 ( .A(n120), .Y(n256) );
  AOI22X1 U308 ( .A0(R1[1]), .A1(n293), .B0(Rin[1]), .B1(n281), .Y(n120) );
  INVX1 U309 ( .A(n121), .Y(n257) );
  AOI22X1 U310 ( .A0(R1[2]), .A1(n292), .B0(Rin[2]), .B1(n282), .Y(n121) );
  INVX1 U311 ( .A(n122), .Y(n258) );
  AOI22X1 U312 ( .A0(R1[3]), .A1(n291), .B0(Rin[3]), .B1(n280), .Y(n122) );
  INVX1 U313 ( .A(n123), .Y(n259) );
  AOI22X1 U314 ( .A0(R1[4]), .A1(n308), .B0(Rin[4]), .B1(n290), .Y(n123) );
  INVX1 U315 ( .A(n124), .Y(n260) );
  AOI22X1 U316 ( .A0(R1[5]), .A1(n297), .B0(Rin[5]), .B1(n280), .Y(n124) );
  INVX1 U317 ( .A(n125), .Y(n261) );
  AOI22X1 U318 ( .A0(R1[6]), .A1(n298), .B0(Rin[6]), .B1(n306), .Y(n125) );
  INVX1 U319 ( .A(n126), .Y(n262) );
  AOI22X1 U320 ( .A0(R1[7]), .A1(n292), .B0(Rin[7]), .B1(n279), .Y(n126) );
  INVX1 U321 ( .A(n127), .Y(n263) );
  AOI22X1 U322 ( .A0(R1[8]), .A1(n302), .B0(Rin[8]), .B1(n285), .Y(n127) );
  INVX1 U323 ( .A(n128), .Y(n264) );
  AOI22X1 U324 ( .A0(R1[9]), .A1(n304), .B0(Rin[9]), .B1(n289), .Y(n128) );
  INVX1 U325 ( .A(n129), .Y(n265) );
  AOI22X1 U326 ( .A0(R1[10]), .A1(n301), .B0(Rin[10]), .B1(n283), .Y(n129) );
  INVX1 U327 ( .A(n130), .Y(n266) );
  AOI22X1 U328 ( .A0(R1[11]), .A1(n295), .B0(Rin[11]), .B1(n279), .Y(n130) );
  INVX1 U329 ( .A(n131), .Y(n267) );
  AOI22X1 U330 ( .A0(R1[12]), .A1(n292), .B0(Rin[12]), .B1(n282), .Y(n131) );
  INVX1 U331 ( .A(n132), .Y(n268) );
  AOI22X1 U332 ( .A0(n272), .A1(n136), .B0(n295), .B1(S2), .Y(n132) );
  AOI22X1 U333 ( .A0(L2[11]), .A1(n300), .B0(l_mux[11]), .B1(n286), .Y(n16) );
endmodule


module mux_13_2to1_3 ( a, b, sel, out );
  input [12:0] a;
  input [12:0] b;
  output [12:0] out;
  input sel;
  wire   n16, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n1,
         n2, n3, n4;

  INVX1 U1 ( .A(n2), .Y(n3) );
  INVX1 U2 ( .A(n1), .Y(n4) );
  INVX1 U3 ( .A(n2), .Y(n1) );
  INVX1 U4 ( .A(sel), .Y(n2) );
  INVX1 U5 ( .A(n29), .Y(out[0]) );
  AOI22X1 U6 ( .A0(a[0]), .A1(n3), .B0(b[0]), .B1(n2), .Y(n29) );
  INVX1 U7 ( .A(n25), .Y(out[1]) );
  AOI22X1 U8 ( .A0(a[1]), .A1(n3), .B0(b[1]), .B1(n2), .Y(n25) );
  INVX1 U9 ( .A(n24), .Y(out[2]) );
  AOI22X1 U10 ( .A0(a[2]), .A1(n3), .B0(b[2]), .B1(n2), .Y(n24) );
  INVX1 U11 ( .A(n23), .Y(out[3]) );
  AOI22X1 U12 ( .A0(a[3]), .A1(n3), .B0(b[3]), .B1(n4), .Y(n23) );
  INVX1 U13 ( .A(n22), .Y(out[4]) );
  AOI22X1 U14 ( .A0(a[4]), .A1(n3), .B0(b[4]), .B1(n4), .Y(n22) );
  INVX1 U15 ( .A(n21), .Y(out[5]) );
  AOI22X1 U16 ( .A0(a[5]), .A1(n3), .B0(b[5]), .B1(n4), .Y(n21) );
  INVX1 U17 ( .A(n20), .Y(out[6]) );
  AOI22X1 U18 ( .A0(a[6]), .A1(n3), .B0(b[6]), .B1(n4), .Y(n20) );
  INVX1 U19 ( .A(n19), .Y(out[7]) );
  AOI22X1 U20 ( .A0(a[7]), .A1(n1), .B0(b[7]), .B1(n2), .Y(n19) );
  INVX1 U21 ( .A(n18), .Y(out[8]) );
  AOI22X1 U22 ( .A0(a[8]), .A1(n1), .B0(b[8]), .B1(n4), .Y(n18) );
  INVX1 U23 ( .A(n16), .Y(out[9]) );
  AOI22X1 U24 ( .A0(sel), .A1(a[9]), .B0(b[9]), .B1(n2), .Y(n16) );
  INVX1 U25 ( .A(n28), .Y(out[10]) );
  AOI22X1 U26 ( .A0(a[10]), .A1(n3), .B0(b[10]), .B1(n4), .Y(n28) );
  INVX1 U27 ( .A(n27), .Y(out[11]) );
  AOI22X1 U28 ( .A0(a[11]), .A1(n3), .B0(b[11]), .B1(n4), .Y(n27) );
  INVX1 U29 ( .A(n26), .Y(out[12]) );
  AOI22X1 U30 ( .A0(a[12]), .A1(n3), .B0(b[12]), .B1(n4), .Y(n26) );
endmodule


module mux_1_2to1_1 ( a, b, sel, out );
  input a, b, sel;
  output out;
  wire   n3;

  OAI2BB2X1 U1 ( .B0(n3), .B1(sel), .A0N(sel), .A1N(a), .Y(out) );
  INVX1 U2 ( .A(b), .Y(n3) );
endmodule


module mux_5_2to1_1 ( a, b, sel, out );
  input [4:0] a;
  input [4:0] b;
  output [4:0] out;
  input sel;
  wire   n8, n10, n11, n12, n13, n1;

  INVX1 U1 ( .A(sel), .Y(n1) );
  INVX1 U2 ( .A(n10), .Y(out[3]) );
  AOI22X1 U3 ( .A0(a[3]), .A1(sel), .B0(b[3]), .B1(n1), .Y(n10) );
  INVX1 U4 ( .A(n11), .Y(out[2]) );
  AOI22X1 U5 ( .A0(a[2]), .A1(sel), .B0(b[2]), .B1(n1), .Y(n11) );
  INVX1 U6 ( .A(n8), .Y(out[4]) );
  AOI22X1 U7 ( .A0(sel), .A1(a[4]), .B0(b[4]), .B1(n1), .Y(n8) );
  INVX1 U8 ( .A(n13), .Y(out[0]) );
  AOI22X1 U9 ( .A0(a[0]), .A1(sel), .B0(b[0]), .B1(n1), .Y(n13) );
  INVX1 U10 ( .A(n12), .Y(out[1]) );
  AOI22X1 U11 ( .A0(a[1]), .A1(sel), .B0(b[1]), .B1(n1), .Y(n12) );
endmodule


module chien_search_p16_t8 ( lambda0, lambda1, lambda2, lambda3, lambda4, 
        lambda5, lambda6, lambda7, lambda8, enable, sigma1, sigma2, sigma3, 
        sigma4, sigma5, sigma6, sigma7, sigma8, sigma9, sigma10, sigma11, 
        sigma12, sigma13, sigma14, sigma15, sigma16, sel, clk, reset );
  input [12:0] lambda0;
  input [12:0] lambda1;
  input [12:0] lambda2;
  input [12:0] lambda3;
  input [12:0] lambda4;
  input [12:0] lambda5;
  input [12:0] lambda6;
  input [12:0] lambda7;
  input [12:0] lambda8;
  output [12:0] sigma1;
  output [12:0] sigma2;
  output [12:0] sigma3;
  output [12:0] sigma4;
  output [12:0] sigma5;
  output [12:0] sigma6;
  output [12:0] sigma7;
  output [12:0] sigma8;
  output [12:0] sigma9;
  output [12:0] sigma10;
  output [12:0] sigma11;
  output [12:0] sigma12;
  output [12:0] sigma13;
  output [12:0] sigma14;
  output [12:0] sigma15;
  output [12:0] sigma16;
  input enable, sel, clk, reset;
  wire   N419, n2, n3, n4, n5, n6, n7, n8, n11, n12, n13, n14, n15, n16, n19,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n43, n44, n45, n46, n51, n52, n53, n54, n55, n56,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n131, n132, n133, n134, n137, n138,
         n139, n140, n141, n142, n145, n146, n147, n148, n149, n150, n151,
         n152, n155, n156, n157, n158, n159, n160, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n219, n220, n221, n222, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n331, n332, n333,
         n334, n335, n336, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n395, n397, n398,
         n399, n400, n401, n402, n403, n405, n406, n407, n408, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n429, n430, n431, n432, n433, n434, n435,
         n437, n438, n439, n440, n443, n445, n446, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n507, n508, n509, n510, n511, n512, n513, n515,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n617, n618, n619, n620, n621, n622, n623, n624,
         n627, n628, n629, n630, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n649, n650, n651, n652,
         n653, n654, n657, n658, n659, n660, n661, n662, n667, n668, n669,
         n670, n673, n674, n675, n676, n677, n678, n681, n682, n683, n684,
         n685, n686, n689, n690, n691, n692, n693, n694, n697, n698, n699,
         n700, n701, n702, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n723, n724, n725, n726, n729,
         n730, n731, n732, n733, n734, n735, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n763, n764, n765,
         n766, n771, n772, n773, n774, n777, n778, n779, n780, n781, n782,
         n785, n786, n787, n788, n789, n790, n791, n793, n794, n795, n796,
         n797, n798, n801, n802, n803, n804, n805, n806, n809, n810, n811,
         n812, n813, n814, n817, n818, n819, n820, n821, n822, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n841, n842, n843, n844, n845, n846, n849, n850, n851, n852,
         n853, n854, n855, n856, n859, n860, n861, n862, n867, n868, n869,
         n870, n873, n874, n875, n876, n877, n878, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n893, n894, n897, n898,
         n899, n900, n901, n902, n905, n906, n907, n908, n909, n910, n911,
         n912, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n930, n931, n932, n933, n934, n937, n938, n939, n940,
         n941, n942, n943, n944, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n968, n971, n972, n973, n974, n975, n976, n978, n979,
         n980, n981, n982, n985, n986, n987, n988, n989, n990, n993, n994,
         n995, n996, n997, n998, n1001, n1002, n1003, n1004, n1005, n1006,
         n1011, n1012, n1013, n1014, n1017, n1018, n1019, n1020, n1021, n1022,
         n1025, n1026, n1027, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1073, n1074, n1075, n1076, n1077, n1078, n1083, n1084, n1085,
         n1086, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1115, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1145, n1146,
         n1147, n1148, n1149, n1150, n1155, n1156, n1157, n1158, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1187, n1188, n1189, n1190, n1193, n1194, n1195, n1196, n1197,
         n1198, n1201, n1202, n1203, n1204, n1205, n1206, n1209, n1210, n1211,
         n1212, n1213, n1214, n1219, n1220, n1221, n1222, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1243, n1244, n1245, n1246, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1267,
         n1268, n1269, n1270, n1273, n1274, n1275, n1276, n1277, n1278, n1281,
         n1282, n1283, n1284, n1285, n1286, n1289, n1290, n1291, n1292, n1293,
         n1294, n1297, n1298, n1299, n1300, n1301, n1302, n1305, n1306, n1307,
         n1308, n1309, n1310, n1313, n1314, n1315, n1316, n1317, n1318, n1321,
         n1322, n1323, n1324, n1325, n1326, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1363, n1364, n1365, n1366, n1367,
         n1368, n1371, n1372, n1373, n1374, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1395,
         n1396, n1397, n1398, n1403, n1404, n1405, n1406, n1409, n1410, n1411,
         n1412, n1413, n1414, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1435, n1436, n1437,
         n1438, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1467, n1468, n1469, n1470, n1471, n1472, n1475, n1476, n1477,
         n1478, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1491,
         n1492, n1493, n1494, n1495, n1496, n1499, n1500, n1501, n1502, n1505,
         n1506, n1507, n1508, n1509, n1510, n1515, n1516, n1517, n1518, n1523,
         n1524, n1525, n1526, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1539, n1540, n1541, n1542, n1547, n1548, n1549, n1550, n1551,
         n1552, n1555, n1556, n1557, n1558, n1559, n1560, n1563, n1564, n1565,
         n1566, n1567, n1568, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1593, n1594, n1595, n1596, n1597, n1598, n1603,
         n1604, n1605, n1606, n1611, n1612, n1613, n1614, n1615, n1616, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1635, n1636, n1637, n1638, n1639, n1640, n1643,
         n1644, n1645, n1646, n1647, n1648, n1651, n1652, n1653, n1654, n1659,
         n1660, n1661, n1662, n1663, n1664, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1, n9, n10, n17, n18, n20, n39, n40, n41, n42,
         n47, n48, n49, n50, n57, n58, n71, n72, n129, n130, n135, n136, n143,
         n144, n153, n154, n161, n162, n193, n194, n217, n218, n223, n224,
         n268, n297, n298, n327, n328, n329, n330, n337, n338, n351, n352,
         n353, n354, n392, n393, n394, n396, n404, n409, n410, n428, n436,
         n441, n442, n444, n447, n448, n463, n464, n476, n489, n490, n505,
         n506, n514, n516, n529, n530, n545, n546, n561, n562, n585, n586,
         n616, n625, n626, n631, n632, n647, n648, n655, n656, n663, n664,
         n665, n666, n671, n672, n679, n680, n687, n688, n695, n696, n703,
         n704, n719, n720, n721, n722, n727, n728, n736, n761, n762, n767,
         n768, n769, n770, n775, n776, n783, n784, n792, n799, n800, n807,
         n808, n815, n816, n823, n824, n839, n840, n847, n848, n857, n858,
         n863, n864, n865, n866, n871, n872, n879, n880, n892, n895, n896,
         n903, n904, n913, n914, n927, n928, n929, n935, n936, n945, n946,
         n967, n969, n970, n977, n983, n984, n991, n992, n999, n1000, n1007,
         n1008, n1009, n1010, n1015, n1016, n1023, n1024, n1028, n1047, n1048,
         n1049, n1050, n1071, n1072, n1079, n1080, n1081, n1082, n1087, n1088,
         n1103, n1104, n1113, n1114, n1116, n1129, n1130, n1143, n1144, n1151,
         n1152, n1153, n1154, n1159, n1160, n1172, n1185, n1186, n1191, n1192,
         n1199, n1200, n1207, n1208, n1215, n1216, n1217, n1218, n1223, n1224,
         n1239, n1240, n1241, n1242, n1247, n1248, n1249, n1250, n1265, n1266,
         n1271, n1272, n1279, n1280, n1287, n1288, n1295, n1296, n1303, n1304,
         n1311, n1312, n1319, n1320, n1327, n1328, n1345, n1346, n1361, n1362,
         n1369, n1370, n1375, n1376, n1391, n1392, n1393, n1394, n1399, n1400,
         n1401, n1402, n1407, n1408, n1415, n1416, n1431, n1432, n1433, n1434,
         n1439, n1440, n1441, n1442, n1455, n1456, n1465, n1466, n1473, n1474,
         n1479, n1480, n1489, n1490, n1497, n1498, n1503, n1504, n1511, n1512,
         n1513, n1514, n1519, n1520, n1521, n1522, n1527, n1528, n1537, n1538,
         n1543, n1544, n1545, n1546, n1553, n1554, n1561, n1562, n1569, n1570,
         n1591, n1592, n1599, n1600, n1601, n1602, n1607, n1608, n1609, n1610,
         n1617, n1618, n1633, n1634, n1641, n1642, n1649, n1650, n1655, n1656,
         n1657, n1658, n1665, n1666, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951;
  wire   [12:0] line1;
  wire   [12:0] line2;
  wire   [12:0] line3;
  wire   [12:0] line4;
  wire   [12:0] line5;
  wire   [12:0] line6;
  wire   [12:0] line7;
  wire   [12:0] line8;
  wire   [12:0] col0;
  wire   [12:0] L16_1;
  wire   [12:0] col1;
  wire   [12:0] L16_2;
  wire   [12:0] col2;
  wire   [12:0] L16_3;
  wire   [12:0] col3;
  wire   [12:0] L16_4;
  wire   [12:0] col4;
  wire   [12:0] L16_5;
  wire   [12:0] col5;
  wire   [12:0] L16_6;
  wire   [12:0] col6;
  wire   [12:0] L16_7;
  wire   [12:0] col7;
  wire   [12:0] L16_8;
  wire   [12:0] col8;
  wire   [12:0] L1_1;
  wire   [12:0] L2_1;
  wire   [12:0] L3_1;
  wire   [12:0] L4_1;
  wire   [12:0] L5_1;
  wire   [12:0] L6_1;
  wire   [12:0] L7_1;
  wire   [12:0] L8_1;
  wire   [12:0] L9_1;
  wire   [12:0] L10_1;
  wire   [12:0] L11_1;
  wire   [12:0] L12_1;
  wire   [12:0] L13_1;
  wire   [12:0] L14_1;
  wire   [12:0] L15_1;
  wire   [12:0] L1_2;
  wire   [12:0] L2_2;
  wire   [12:0] L3_2;
  wire   [12:0] L4_2;
  wire   [12:0] L5_2;
  wire   [12:0] L6_2;
  wire   [12:0] L7_2;
  wire   [12:0] L8_2;
  wire   [12:0] L9_2;
  wire   [12:0] L10_2;
  wire   [12:0] L11_2;
  wire   [12:0] L12_2;
  wire   [12:0] L13_2;
  wire   [12:0] L14_2;
  wire   [12:0] L15_2;
  wire   [12:0] L1_3;
  wire   [12:0] L2_3;
  wire   [12:0] L3_3;
  wire   [12:0] L4_3;
  wire   [12:0] L5_3;
  wire   [12:0] L6_3;
  wire   [12:0] L7_3;
  wire   [12:0] L8_3;
  wire   [12:0] L9_3;
  wire   [12:0] L10_3;
  wire   [12:0] L11_3;
  wire   [12:0] L12_3;
  wire   [12:0] L13_3;
  wire   [12:0] L14_3;
  wire   [12:0] L15_3;
  wire   [12:0] L1_4;
  wire   [12:0] L2_4;
  wire   [12:0] L3_4;
  wire   [12:0] L4_4;
  wire   [12:0] L5_4;
  wire   [12:0] L6_4;
  wire   [12:0] L7_4;
  wire   [12:0] L8_4;
  wire   [12:0] L9_4;
  wire   [12:0] L10_4;
  wire   [12:0] L11_4;
  wire   [12:0] L12_4;
  wire   [12:0] L13_4;
  wire   [12:0] L14_4;
  wire   [12:0] L15_4;
  wire   [12:0] L1_5;
  wire   [12:0] L2_5;
  wire   [12:0] L3_5;
  wire   [12:0] L4_5;
  wire   [12:0] L5_5;
  wire   [12:0] L6_5;
  wire   [12:0] L7_5;
  wire   [12:0] L8_5;
  wire   [12:0] L9_5;
  wire   [12:0] L10_5;
  wire   [12:0] L11_5;
  wire   [12:0] L12_5;
  wire   [12:0] L13_5;
  wire   [12:0] L14_5;
  wire   [12:0] L15_5;
  wire   [12:0] L1_6;
  wire   [12:0] L2_6;
  wire   [12:0] L3_6;
  wire   [12:0] L4_6;
  wire   [12:0] L5_6;
  wire   [12:0] L6_6;
  wire   [12:0] L7_6;
  wire   [12:0] L8_6;
  wire   [12:0] L9_6;
  wire   [12:0] L10_6;
  wire   [12:0] L11_6;
  wire   [12:0] L12_6;
  wire   [12:0] L13_6;
  wire   [12:0] L14_6;
  wire   [12:0] L15_6;
  wire   [12:0] L1_7;
  wire   [12:0] L2_7;
  wire   [12:0] L3_7;
  wire   [12:0] L4_7;
  wire   [12:0] L5_7;
  wire   [12:0] L6_7;
  wire   [12:0] L7_7;
  wire   [12:0] L8_7;
  wire   [12:0] L9_7;
  wire   [12:0] L10_7;
  wire   [12:0] L11_7;
  wire   [12:0] L12_7;
  wire   [12:0] L13_7;
  wire   [12:0] L14_7;
  wire   [12:0] L15_7;
  wire   [12:0] L1_8;
  wire   [12:0] L2_8;
  wire   [12:0] L3_8;
  wire   [12:0] L4_8;
  wire   [12:0] L5_8;
  wire   [12:0] L6_8;
  wire   [12:0] L7_8;
  wire   [12:0] L8_8;
  wire   [12:0] L9_8;
  wire   [12:0] L10_8;
  wire   [12:0] L11_8;
  wire   [12:0] L12_8;
  wire   [12:0] L13_8;
  wire   [12:0] L14_8;
  wire   [12:0] L15_8;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign N419 = enable;

  DFFRHQX4 \sigma16_reg[0]  ( .D(n1823), .CK(clk), .RN(reset), .Q(sigma16[0])
         );
  DFFRHQX4 \sigma9_reg[10]  ( .D(n1716), .CK(clk), .RN(reset), .Q(sigma9[10])
         );
  XNOR2X4 U592 ( .A(L16_2[0]), .B(n1), .Y(n528) );
  multiply_3967 m1 ( .a(lambda1), .c(line1) );
  multiply_7934 m2 ( .a(lambda2), .c(line2) );
  multiply_3710 m3 ( .a(lambda3), .c(line3) );
  multiply_7677 m4 ( .a(lambda4), .c(line4) );
  multiply_3453 m5 ( .a(lambda5), .c(line5) );
  multiply_7420 m6 ( .a(lambda6), .c(line6) );
  multiply_3196 m7 ( .a(lambda7), .c(line7) );
  multiply_7163 m8 ( .a(lambda8), .c(line8) );
  mux13_13_8 mmm0 ( .a(lambda0), .b({n41, n143, n135, n57, n161, n49, n39, n47, 
        n153, n129, n71, n18, n193}), .sel(n10), .enable(N419), .out(col0), 
        .clk(clk), .reset(reset) );
  mux13_13_7 mmm1 ( .a(line1), .b({L16_1[12:1], n1}), .sel(n10), .enable(N419), 
        .out(col1), .clk(clk), .reset(reset) );
  mux13_13_6 mmm2 ( .a(line2), .b(L16_2), .sel(n10), .enable(N419), .out(col2), 
        .clk(clk), .reset(reset) );
  mux13_13_5 mmm3 ( .a(line3), .b(L16_3), .sel(sel), .enable(N419), .out(col3), 
        .clk(clk), .reset(reset) );
  mux13_13_4 mmm4 ( .a(line4), .b(L16_4), .sel(sel), .enable(N419), .out(col4), 
        .clk(clk), .reset(reset) );
  mux13_13_3 mmm5 ( .a(line5), .b(L16_5), .sel(n10), .enable(N419), .out(col5), 
        .clk(clk), .reset(reset) );
  mux13_13_2 mmm6 ( .a(line6), .b(L16_6), .sel(n10), .enable(N419), .out(col6), 
        .clk(clk), .reset(reset) );
  mux13_13_1 mmm7 ( .a(line7), .b({L16_7[12:3], n1903, L16_7[1:0]}), .sel(sel), 
        .enable(N419), .out(col7), .clk(clk), .reset(reset) );
  mux13_13_0 mmm8 ( .a(line8), .b(L16_8), .sel(sel), .enable(N419), .out(col8), 
        .clk(clk), .reset(reset) );
  multiplier_column1_p16 c1 ( .b(col1), .P1({L1_1[12:10], 
        SYNOPSYS_UNCONNECTED__0, L1_1[8:0]}), .P2(L2_1), .P3(L3_1), .P4(L4_1), 
        .P5(L5_1), .P6(L6_1), .P7(L7_1), .P8(L8_1), .P9(L9_1), .P10(L10_1), 
        .P11(L11_1), .P12(L12_1), .P13(L13_1), .P14(L14_1), .P15(L15_1), .P16(
        L16_1) );
  multiplier_column2_p16 c2 ( .b(col2), .P1(L1_2), .P2(L2_2), .P3(L3_2), .P4({
        SYNOPSYS_UNCONNECTED__1, L4_2[11:0]}), .P5(L5_2), .P6(L6_2), .P7(L7_2), 
        .P8(L8_2), .P9(L9_2), .P10(L10_2), .P11(L11_2), .P12(L12_2), .P13(
        L13_2), .P14(L14_2), .P15(L15_2), .P16(L16_2) );
  multiplier_column3_p16 c3 ( .b(col3), .P1(L1_3), .P2(L2_3), .P3(L3_3), .P4(
        L4_3), .P5(L5_3), .P6(L6_3), .P7(L7_3), .P8(L8_3), .P9(L9_3), .P10(
        L10_3), .P11(L11_3), .P12(L12_3), .P13(L13_3), .P14(L14_3), .P15(L15_3), .P16(L16_3) );
  multiplier_column4_p16 c4 ( .b(col4), .P1(L1_4), .P2(L2_4), .P3(L3_4), .P4(
        L4_4), .P5(L5_4), .P6(L6_4), .P7(L7_4), .P8(L8_4), .P9(L9_4), .P10(
        L10_4), .P11(L11_4), .P12(L12_4), .P13(L13_4), .P14(L14_4), .P15(L15_4), .P16(L16_4) );
  multiplier_column5_p16 c5 ( .b(col5), .P1(L1_5), .P2(L2_5), .P3(L3_5), .P4(
        L4_5), .P5(L5_5), .P6(L6_5), .P7(L7_5), .P8(L8_5), .P9(L9_5), .P10(
        L10_5), .P11(L11_5), .P12(L12_5), .P13(L13_5), .P14(L14_5), .P15(L15_5), .P16(L16_5) );
  multiplier_column6_p16 c6 ( .b(col6), .P1(L1_6), .P2(L2_6), .P3(L3_6), .P4(
        L4_6), .P5(L5_6), .P6(L6_6), .P7(L7_6), .P8(L8_6), .P9(L9_6), .P10(
        L10_6), .P11(L11_6), .P12(L12_6), .P13(L13_6), .P14(L14_6), .P15(L15_6), .P16(L16_6) );
  multiplier_column7_p16 c7 ( .b({col7[12:9], n1904, col7[7:0]}), .P1(L1_7), 
        .P2(L2_7), .P3(L3_7), .P4(L4_7), .P5(L5_7), .P6(L6_7), .P7(L7_7), .P8(
        L8_7), .P9(L9_7), .P10(L10_7), .P11(L11_7), .P12(L12_7), .P13(L13_7), 
        .P14(L14_7), .P15(L15_7), .P16(L16_7) );
  multiplier_column8_p16 c8 ( .b(col8), .P1(L1_8), .P2(L2_8), .P3(L3_8), .P4(
        L4_8), .P5(L5_8), .P6(L6_8), .P7(L7_8), .P8(L8_8), .P9(L9_8), .P10(
        L10_8), .P11(L11_8), .P12(L12_8), .P13(L13_8), .P14(L14_8), .P15(L15_8), .P16(L16_8) );
  DFFRHQX1 \sigma6_reg[12]  ( .D(n1757), .CK(clk), .RN(reset), .Q(sigma6[12])
         );
  DFFRHQX1 \sigma4_reg[1]  ( .D(n1772), .CK(clk), .RN(reset), .Q(sigma4[1]) );
  DFFRHQX1 \sigma6_reg[2]  ( .D(n1747), .CK(clk), .RN(reset), .Q(sigma6[2]) );
  DFFRHQX1 \sigma10_reg[12]  ( .D(n1705), .CK(clk), .RN(reset), .Q(sigma10[12]) );
  DFFRHQX1 \sigma16_reg[9]  ( .D(n1832), .CK(clk), .RN(reset), .Q(sigma16[9])
         );
  DFFRHQX1 \sigma16_reg[6]  ( .D(n1829), .CK(clk), .RN(reset), .Q(sigma16[6])
         );
  DFFRHQX1 \sigma4_reg[4]  ( .D(n1775), .CK(clk), .RN(reset), .Q(sigma4[4]) );
  DFFRHQX1 \sigma3_reg[11]  ( .D(n1795), .CK(clk), .RN(reset), .Q(sigma3[11])
         );
  DFFRHQX1 \sigma3_reg[8]  ( .D(n1792), .CK(clk), .RN(reset), .Q(sigma3[8]) );
  DFFRHQX1 \sigma4_reg[11]  ( .D(n1782), .CK(clk), .RN(reset), .Q(sigma4[11])
         );
  DFFRHQX1 \sigma4_reg[8]  ( .D(n1779), .CK(clk), .RN(reset), .Q(sigma4[8]) );
  DFFRHQX1 \sigma10_reg[11]  ( .D(n1704), .CK(clk), .RN(reset), .Q(sigma10[11]) );
  DFFRHQX1 \sigma2_reg[12]  ( .D(n1809), .CK(clk), .RN(reset), .Q(sigma2[12])
         );
  DFFRHQX1 \sigma3_reg[7]  ( .D(n1791), .CK(clk), .RN(reset), .Q(sigma3[7]) );
  DFFRHQX1 \sigma4_reg[10]  ( .D(n1781), .CK(clk), .RN(reset), .Q(sigma4[10])
         );
  DFFRHQX1 \sigma4_reg[7]  ( .D(n1778), .CK(clk), .RN(reset), .Q(sigma4[7]) );
  DFFRHQX1 \sigma5_reg[4]  ( .D(n1762), .CK(clk), .RN(reset), .Q(sigma5[4]) );
  DFFRHQX1 \sigma8_reg[10]  ( .D(n1729), .CK(clk), .RN(reset), .Q(sigma8[10])
         );
  DFFRHQX1 \sigma8_reg[7]  ( .D(n1726), .CK(clk), .RN(reset), .Q(sigma8[7]) );
  DFFRHQX1 \sigma10_reg[10]  ( .D(n1703), .CK(clk), .RN(reset), .Q(sigma10[10]) );
  DFFRHQX1 \sigma10_reg[7]  ( .D(n1700), .CK(clk), .RN(reset), .Q(sigma10[7])
         );
  DFFRHQX1 \sigma10_reg[4]  ( .D(n1697), .CK(clk), .RN(reset), .Q(sigma10[4])
         );
  DFFRHQX1 \sigma2_reg[1]  ( .D(n1798), .CK(clk), .RN(reset), .Q(sigma2[1]) );
  DFFRHQX1 \sigma13_reg[8]  ( .D(n1870), .CK(clk), .RN(reset), .Q(sigma13[8])
         );
  DFFRHQX1 \sigma13_reg[5]  ( .D(n1867), .CK(clk), .RN(reset), .Q(sigma13[5])
         );
  DFFRHQX1 \sigma13_reg[3]  ( .D(n1865), .CK(clk), .RN(reset), .Q(sigma13[3])
         );
  DFFRHQX1 \sigma16_reg[12]  ( .D(n1835), .CK(clk), .RN(reset), .Q(sigma16[12]) );
  DFFRHQX1 \sigma16_reg[8]  ( .D(n1831), .CK(clk), .RN(reset), .Q(sigma16[8])
         );
  DFFRHQX1 \sigma16_reg[3]  ( .D(n1826), .CK(clk), .RN(reset), .Q(sigma16[3])
         );
  DFFRHQX1 \sigma2_reg[4]  ( .D(n1801), .CK(clk), .RN(reset), .Q(sigma2[4]) );
  DFFRHQX1 \sigma3_reg[3]  ( .D(n1787), .CK(clk), .RN(reset), .Q(sigma3[3]) );
  DFFRHQX1 \sigma4_reg[5]  ( .D(n1776), .CK(clk), .RN(reset), .Q(sigma4[5]) );
  DFFRHQX1 \sigma4_reg[3]  ( .D(n1774), .CK(clk), .RN(reset), .Q(sigma4[3]) );
  DFFRHQX1 \sigma7_reg[5]  ( .D(n1737), .CK(clk), .RN(reset), .Q(sigma7[5]) );
  DFFRHQX1 \sigma7_reg[1]  ( .D(n1733), .CK(clk), .RN(reset), .Q(sigma7[1]) );
  DFFRHQX1 \sigma8_reg[5]  ( .D(n1724), .CK(clk), .RN(reset), .Q(sigma8[5]) );
  DFFRHQX1 \sigma8_reg[1]  ( .D(n1720), .CK(clk), .RN(reset), .Q(sigma8[1]) );
  DFFRHQX1 \sigma12_reg[12]  ( .D(n1679), .CK(clk), .RN(reset), .Q(sigma12[12]) );
  DFFRHQX1 \sigma12_reg[3]  ( .D(n1670), .CK(clk), .RN(reset), .Q(sigma12[3])
         );
  DFFRHQX1 \sigma1_reg[9]  ( .D(n1819), .CK(clk), .RN(reset), .Q(sigma1[9]) );
  DFFRHQX1 \sigma1_reg[6]  ( .D(n1816), .CK(clk), .RN(reset), .Q(sigma1[6]) );
  DFFRHQX1 \sigma2_reg[11]  ( .D(n1808), .CK(clk), .RN(reset), .Q(sigma2[11])
         );
  DFFRHQX1 \sigma2_reg[8]  ( .D(n1805), .CK(clk), .RN(reset), .Q(sigma2[8]) );
  DFFRHQX1 \sigma3_reg[12]  ( .D(n1796), .CK(clk), .RN(reset), .Q(sigma3[12])
         );
  DFFRHQX1 \sigma3_reg[9]  ( .D(n1793), .CK(clk), .RN(reset), .Q(sigma3[9]) );
  DFFRHQX1 \sigma4_reg[12]  ( .D(n1783), .CK(clk), .RN(reset), .Q(sigma4[12])
         );
  DFFRHQX1 \sigma4_reg[9]  ( .D(n1780), .CK(clk), .RN(reset), .Q(sigma4[9]) );
  DFFRHQX1 \sigma5_reg[9]  ( .D(n1767), .CK(clk), .RN(reset), .Q(sigma5[9]) );
  DFFRHQX1 \sigma7_reg[12]  ( .D(n1744), .CK(clk), .RN(reset), .Q(sigma7[12])
         );
  DFFRHQX1 \sigma8_reg[12]  ( .D(n1731), .CK(clk), .RN(reset), .Q(sigma8[12])
         );
  DFFRHQX1 \sigma8_reg[9]  ( .D(n1728), .CK(clk), .RN(reset), .Q(sigma8[9]) );
  DFFRHQX1 \sigma10_reg[9]  ( .D(n1702), .CK(clk), .RN(reset), .Q(sigma10[9])
         );
  DFFRHQX1 \sigma10_reg[6]  ( .D(n1699), .CK(clk), .RN(reset), .Q(sigma10[6])
         );
  DFFRHQX1 \sigma2_reg[2]  ( .D(n1799), .CK(clk), .RN(reset), .Q(sigma2[2]) );
  DFFRHQX1 \sigma2_reg[0]  ( .D(n1797), .CK(clk), .RN(reset), .Q(sigma2[0]) );
  DFFRHQX1 \sigma3_reg[0]  ( .D(n1784), .CK(clk), .RN(reset), .Q(sigma3[0]) );
  DFFRHQX1 \sigma12_reg[1]  ( .D(n1668), .CK(clk), .RN(reset), .Q(sigma12[1])
         );
  DFFRHQX1 \sigma13_reg[6]  ( .D(n1868), .CK(clk), .RN(reset), .Q(sigma13[6])
         );
  DFFRHQX1 \sigma13_reg[1]  ( .D(n1863), .CK(clk), .RN(reset), .Q(sigma13[1])
         );
  DFFRHQX1 \sigma3_reg[4]  ( .D(n1788), .CK(clk), .RN(reset), .Q(sigma3[4]) );
  DFFRHQX1 \sigma3_reg[2]  ( .D(n1786), .CK(clk), .RN(reset), .Q(sigma3[2]) );
  DFFRHQX1 \sigma4_reg[2]  ( .D(n1773), .CK(clk), .RN(reset), .Q(sigma4[2]) );
  DFFRHQX1 \sigma4_reg[0]  ( .D(n1771), .CK(clk), .RN(reset), .Q(sigma4[0]) );
  DFFRHQX1 \sigma7_reg[2]  ( .D(n1734), .CK(clk), .RN(reset), .Q(sigma7[2]) );
  DFFRHQX1 \sigma7_reg[0]  ( .D(n1732), .CK(clk), .RN(reset), .Q(sigma7[0]) );
  DFFRHQX1 \sigma8_reg[2]  ( .D(n1721), .CK(clk), .RN(reset), .Q(sigma8[2]) );
  DFFRHQX1 \sigma12_reg[9]  ( .D(n1676), .CK(clk), .RN(reset), .Q(sigma12[9])
         );
  DFFRHQX1 \sigma16_reg[2]  ( .D(n1825), .CK(clk), .RN(reset), .Q(sigma16[2])
         );
  DFFRHQX1 \sigma1_reg[2]  ( .D(n1812), .CK(clk), .RN(reset), .Q(sigma1[2]) );
  DFFRHQX1 \sigma5_reg[2]  ( .D(n1760), .CK(clk), .RN(reset), .Q(sigma5[2]) );
  DFFRHQX1 \sigma10_reg[2]  ( .D(n1695), .CK(clk), .RN(reset), .Q(sigma10[2])
         );
  DFFRHQX1 \sigma10_reg[3]  ( .D(n1696), .CK(clk), .RN(reset), .Q(sigma10[3])
         );
  DFFRHQX1 \sigma12_reg[0]  ( .D(n1667), .CK(clk), .RN(reset), .Q(sigma12[0])
         );
  DFFRHQX1 \sigma11_reg[10]  ( .D(n1690), .CK(clk), .RN(reset), .Q(sigma11[10]) );
  DFFRHQX1 \sigma13_reg[7]  ( .D(n1869), .CK(clk), .RN(reset), .Q(sigma13[7])
         );
  DFFRHQX1 \sigma13_reg[2]  ( .D(n1864), .CK(clk), .RN(reset), .Q(sigma13[2])
         );
  DFFRHQX1 \sigma2_reg[5]  ( .D(n1802), .CK(clk), .RN(reset), .Q(sigma2[5]) );
  DFFRHQX1 \sigma4_reg[6]  ( .D(n1777), .CK(clk), .RN(reset), .Q(sigma4[6]) );
  DFFRHQX1 \sigma7_reg[6]  ( .D(n1738), .CK(clk), .RN(reset), .Q(sigma7[6]) );
  DFFRHQX1 \sigma8_reg[6]  ( .D(n1725), .CK(clk), .RN(reset), .Q(sigma8[6]) );
  DFFRHQX1 \sigma12_reg[2]  ( .D(n1669), .CK(clk), .RN(reset), .Q(sigma12[2])
         );
  DFFRHQX1 \sigma11_reg[0]  ( .D(n1680), .CK(clk), .RN(reset), .Q(sigma11[0])
         );
  DFFRHQX1 \sigma15_reg[7]  ( .D(n1856), .CK(clk), .RN(reset), .Q(sigma15[7])
         );
  DFFRHQX1 \sigma15_reg[6]  ( .D(n1855), .CK(clk), .RN(reset), .Q(sigma15[6])
         );
  DFFRHQX1 \sigma14_reg[8]  ( .D(n1844), .CK(clk), .RN(reset), .Q(sigma14[8])
         );
  DFFRHQX1 \sigma14_reg[7]  ( .D(n1843), .CK(clk), .RN(reset), .Q(sigma14[7])
         );
  DFFRHQX1 \sigma14_reg[3]  ( .D(n1839), .CK(clk), .RN(reset), .Q(sigma14[3])
         );
  DFFRHQX1 \sigma15_reg[9]  ( .D(n1858), .CK(clk), .RN(reset), .Q(sigma15[9])
         );
  DFFRHQX1 \sigma15_reg[2]  ( .D(n1851), .CK(clk), .RN(reset), .Q(sigma15[2])
         );
  DFFRHQX1 \sigma13_reg[11]  ( .D(n1873), .CK(clk), .RN(reset), .Q(sigma13[11]) );
  DFFRHQX1 \sigma11_reg[11]  ( .D(n1691), .CK(clk), .RN(reset), .Q(sigma11[11]) );
  DFFRHQX1 \sigma3_reg[6]  ( .D(n1790), .CK(clk), .RN(reset), .Q(sigma3[6]) );
  DFFRHQX1 \sigma2_reg[3]  ( .D(n1800), .CK(clk), .RN(reset), .Q(sigma2[3]) );
  DFFRHQX1 \sigma3_reg[1]  ( .D(n1785), .CK(clk), .RN(reset), .Q(sigma3[1]) );
  DFFRHQX1 \sigma3_reg[10]  ( .D(n1794), .CK(clk), .RN(reset), .Q(sigma3[10])
         );
  DFFRHQX2 \sigma1_reg[0]  ( .D(n1810), .CK(clk), .RN(reset), .Q(sigma1[0]) );
  DFFRHQX4 \sigma7_reg[11]  ( .D(n1743), .CK(clk), .RN(reset), .Q(sigma7[11])
         );
  DFFRHQX4 \sigma6_reg[9]  ( .D(n1754), .CK(clk), .RN(reset), .Q(sigma6[9]) );
  DFFRHQX2 \sigma6_reg[1]  ( .D(n1746), .CK(clk), .RN(reset), .Q(sigma6[1]) );
  DFFRHQX1 \sigma16_reg[5]  ( .D(n1828), .CK(clk), .RN(reset), .Q(sigma16[5])
         );
  DFFRHQX4 \sigma6_reg[7]  ( .D(n1752), .CK(clk), .RN(reset), .Q(sigma6[7]) );
  DFFRHQX4 \sigma8_reg[8]  ( .D(n1727), .CK(clk), .RN(reset), .Q(sigma8[8]) );
  DFFRHQX4 \sigma9_reg[11]  ( .D(n1717), .CK(clk), .RN(reset), .Q(sigma9[11])
         );
  DFFRHQX4 \sigma9_reg[12]  ( .D(n1718), .CK(clk), .RN(reset), .Q(sigma9[12])
         );
  DFFRHQX4 \sigma9_reg[9]  ( .D(n1715), .CK(clk), .RN(reset), .Q(sigma9[9]) );
  DFFRHQX4 \sigma11_reg[5]  ( .D(n1685), .CK(clk), .RN(reset), .Q(sigma11[5])
         );
  DFFRHQX4 \sigma16_reg[11]  ( .D(n1834), .CK(clk), .RN(reset), .Q(sigma16[11]) );
  DFFRHQX4 \sigma5_reg[8]  ( .D(n1766), .CK(clk), .RN(reset), .Q(sigma5[8]) );
  DFFRHQX2 \sigma1_reg[11]  ( .D(n1821), .CK(clk), .RN(reset), .Q(sigma1[11])
         );
  DFFRHQX4 \sigma13_reg[12]  ( .D(n1874), .CK(clk), .RN(reset), .Q(sigma13[12]) );
  DFFRHQX4 \sigma6_reg[8]  ( .D(n1753), .CK(clk), .RN(reset), .Q(sigma6[8]) );
  DFFRHQX4 \sigma5_reg[1]  ( .D(n1759), .CK(clk), .RN(reset), .Q(sigma5[1]) );
  DFFRHQX4 \sigma11_reg[4]  ( .D(n1684), .CK(clk), .RN(reset), .Q(sigma11[4])
         );
  DFFRHQX4 \sigma5_reg[6]  ( .D(n1764), .CK(clk), .RN(reset), .Q(sigma5[6]) );
  DFFRHQX2 \sigma10_reg[1]  ( .D(n1694), .CK(clk), .RN(reset), .Q(sigma10[1])
         );
  DFFRHQX4 \sigma11_reg[3]  ( .D(n1683), .CK(clk), .RN(reset), .Q(sigma11[3])
         );
  DFFRHQX2 \sigma1_reg[10]  ( .D(n1820), .CK(clk), .RN(reset), .Q(sigma1[10])
         );
  DFFRHQX4 \sigma14_reg[2]  ( .D(n1838), .CK(clk), .RN(reset), .Q(sigma14[2])
         );
  DFFRHQX4 \sigma15_reg[3]  ( .D(n1852), .CK(clk), .RN(reset), .Q(sigma15[3])
         );
  DFFRHQX4 \sigma6_reg[11]  ( .D(n1756), .CK(clk), .RN(reset), .Q(sigma6[11])
         );
  DFFRHQX2 \sigma9_reg[0]  ( .D(n1706), .CK(clk), .RN(reset), .Q(sigma9[0]) );
  DFFRHQX2 \sigma2_reg[7]  ( .D(n1804), .CK(clk), .RN(reset), .Q(sigma2[7]) );
  DFFRHQX4 \sigma16_reg[10]  ( .D(n1833), .CK(clk), .RN(reset), .Q(sigma16[10]) );
  DFFRHQX2 \sigma2_reg[10]  ( .D(n1807), .CK(clk), .RN(reset), .Q(sigma2[10])
         );
  DFFRHQX2 \sigma1_reg[3]  ( .D(n1813), .CK(clk), .RN(reset), .Q(sigma1[3]) );
  DFFRHQX2 \sigma2_reg[9]  ( .D(n1806), .CK(clk), .RN(reset), .Q(sigma2[9]) );
  DFFRHQX4 \sigma1_reg[1]  ( .D(n1811), .CK(clk), .RN(reset), .Q(sigma1[1]) );
  DFFRHQX4 \sigma8_reg[11]  ( .D(n1730), .CK(clk), .RN(reset), .Q(sigma8[11])
         );
  DFFRHQX4 \sigma13_reg[10]  ( .D(n1872), .CK(clk), .RN(reset), .Q(sigma13[10]) );
  DFFRHQX2 \sigma11_reg[6]  ( .D(n1686), .CK(clk), .RN(reset), .Q(sigma11[6])
         );
  DFFRHQX2 \sigma1_reg[4]  ( .D(n1814), .CK(clk), .RN(reset), .Q(sigma1[4]) );
  DFFRHQX1 \sigma7_reg[4]  ( .D(n1736), .CK(clk), .RN(reset), .Q(sigma7[4]) );
  DFFRHQX2 \sigma15_reg[12]  ( .D(n1861), .CK(clk), .RN(reset), .Q(sigma15[12]) );
  DFFRHQX2 \sigma15_reg[4]  ( .D(n1853), .CK(clk), .RN(reset), .Q(sigma15[4])
         );
  DFFRHQX2 \sigma15_reg[11]  ( .D(n1860), .CK(clk), .RN(reset), .Q(sigma15[11]) );
  DFFRHQX2 \sigma14_reg[1]  ( .D(n1837), .CK(clk), .RN(reset), .Q(sigma14[1])
         );
  DFFRHQX2 \sigma11_reg[12]  ( .D(n1692), .CK(clk), .RN(reset), .Q(sigma11[12]) );
  DFFRHQX2 \sigma6_reg[0]  ( .D(n1745), .CK(clk), .RN(reset), .Q(sigma6[0]) );
  DFFRHQX2 \sigma6_reg[5]  ( .D(n1750), .CK(clk), .RN(reset), .Q(sigma6[5]) );
  DFFRHQX1 \sigma13_reg[0]  ( .D(n1862), .CK(clk), .RN(reset), .Q(sigma13[0])
         );
  DFFRHQX2 \sigma11_reg[1]  ( .D(n1681), .CK(clk), .RN(reset), .Q(sigma11[1])
         );
  DFFRHQX2 \sigma1_reg[8]  ( .D(n1818), .CK(clk), .RN(reset), .Q(sigma1[8]) );
  DFFRHQX2 \sigma11_reg[8]  ( .D(n1688), .CK(clk), .RN(reset), .Q(sigma11[8])
         );
  DFFRHQX2 \sigma9_reg[2]  ( .D(n1708), .CK(clk), .RN(reset), .Q(sigma9[2]) );
  DFFRHQX1 \sigma14_reg[4]  ( .D(n1840), .CK(clk), .RN(reset), .Q(sigma14[4])
         );
  DFFRHQX1 \sigma2_reg[6]  ( .D(n1803), .CK(clk), .RN(reset), .Q(sigma2[6]) );
  DFFRHQX2 \sigma9_reg[5]  ( .D(n1711), .CK(clk), .RN(reset), .Q(sigma9[5]) );
  DFFRHQX1 \sigma16_reg[1]  ( .D(n1824), .CK(clk), .RN(reset), .Q(sigma16[1])
         );
  DFFRHQX2 \sigma11_reg[2]  ( .D(n1682), .CK(clk), .RN(reset), .Q(sigma11[2])
         );
  DFFRHQX1 \sigma7_reg[3]  ( .D(n1735), .CK(clk), .RN(reset), .Q(sigma7[3]) );
  DFFRHQX2 \sigma9_reg[3]  ( .D(n1709), .CK(clk), .RN(reset), .Q(sigma9[3]) );
  DFFRHQX1 \sigma12_reg[10]  ( .D(n1677), .CK(clk), .RN(reset), .Q(sigma12[10]) );
  DFFRHQX1 \sigma5_reg[12]  ( .D(n1770), .CK(clk), .RN(reset), .Q(sigma5[12])
         );
  DFFRHQX1 \sigma10_reg[8]  ( .D(n1701), .CK(clk), .RN(reset), .Q(sigma10[8])
         );
  DFFRHQX1 \sigma12_reg[7]  ( .D(n1674), .CK(clk), .RN(reset), .Q(sigma12[7])
         );
  DFFRHQXL \sigma16_reg[7]  ( .D(n1830), .CK(clk), .RN(reset), .Q(sigma16[7])
         );
  DFFRHQX1 \sigma9_reg[7]  ( .D(n1713), .CK(clk), .RN(reset), .Q(sigma9[7]) );
  DFFRHQX1 \sigma5_reg[5]  ( .D(n1763), .CK(clk), .RN(reset), .Q(sigma5[5]) );
  DFFRHQX1 \sigma9_reg[6]  ( .D(n1712), .CK(clk), .RN(reset), .Q(sigma9[6]) );
  DFFRHQX1 \sigma7_reg[7]  ( .D(n1739), .CK(clk), .RN(reset), .Q(sigma7[7]) );
  DFFRHQX1 \sigma14_reg[9]  ( .D(n1845), .CK(clk), .RN(reset), .Q(sigma14[9])
         );
  DFFRHQX1 \sigma12_reg[8]  ( .D(n1675), .CK(clk), .RN(reset), .Q(sigma12[8])
         );
  DFFRHQX1 \sigma9_reg[4]  ( .D(n1710), .CK(clk), .RN(reset), .Q(sigma9[4]) );
  DFFRHQX2 \sigma14_reg[11]  ( .D(n1847), .CK(clk), .RN(reset), .Q(sigma14[11]) );
  DFFRHQX4 \sigma6_reg[10]  ( .D(n1755), .CK(clk), .RN(reset), .Q(sigma6[10])
         );
  DFFRHQX4 \sigma7_reg[8]  ( .D(n1740), .CK(clk), .RN(reset), .Q(sigma7[8]) );
  DFFRHQX4 \sigma13_reg[9]  ( .D(n1871), .CK(clk), .RN(reset), .Q(sigma13[9])
         );
  DFFRHQX4 \sigma8_reg[4]  ( .D(n1723), .CK(clk), .RN(reset), .Q(sigma8[4]) );
  DFFRHQX4 \sigma9_reg[8]  ( .D(n1714), .CK(clk), .RN(reset), .Q(sigma9[8]) );
  DFFRHQX1 \sigma16_reg[4]  ( .D(n1827), .CK(clk), .RN(reset), .Q(sigma16[4])
         );
  DFFRHQX1 \sigma6_reg[6]  ( .D(n1751), .CK(clk), .RN(reset), .Q(sigma6[6]) );
  DFFRHQX2 \sigma15_reg[10]  ( .D(n1859), .CK(clk), .RN(reset), .Q(sigma15[10]) );
  DFFRHQX2 \sigma11_reg[9]  ( .D(n1689), .CK(clk), .RN(reset), .Q(sigma11[9])
         );
  DFFRHQX1 \sigma12_reg[4]  ( .D(n1671), .CK(clk), .RN(reset), .Q(sigma12[4])
         );
  DFFRHQX1 \sigma5_reg[7]  ( .D(n1765), .CK(clk), .RN(reset), .Q(sigma5[7]) );
  DFFRHQX1 \sigma6_reg[3]  ( .D(n1748), .CK(clk), .RN(reset), .Q(sigma6[3]) );
  DFFRHQX1 \sigma10_reg[5]  ( .D(n1698), .CK(clk), .RN(reset), .Q(sigma10[5])
         );
  DFFRHQX1 \sigma3_reg[5]  ( .D(n1789), .CK(clk), .RN(reset), .Q(sigma3[5]) );
  DFFRHQX4 \sigma12_reg[11]  ( .D(n1678), .CK(clk), .RN(reset), .Q(sigma12[11]) );
  DFFRHQX4 \sigma14_reg[12]  ( .D(n1848), .CK(clk), .RN(reset), .Q(sigma14[12]) );
  DFFRHQX4 \sigma12_reg[6]  ( .D(n1673), .CK(clk), .RN(reset), .Q(sigma12[6])
         );
  DFFRHQX4 \sigma6_reg[4]  ( .D(n1749), .CK(clk), .RN(reset), .Q(sigma6[4]) );
  DFFRHQX4 \sigma8_reg[0]  ( .D(n1719), .CK(clk), .RN(reset), .Q(sigma8[0]) );
  DFFRHQX1 \sigma15_reg[0]  ( .D(n1849), .CK(clk), .RN(reset), .Q(sigma15[0])
         );
  DFFRHQX2 \sigma14_reg[5]  ( .D(n1841), .CK(clk), .RN(reset), .Q(sigma14[5])
         );
  DFFRHQX2 \sigma1_reg[5]  ( .D(n1815), .CK(clk), .RN(reset), .Q(sigma1[5]) );
  DFFRHQX1 \sigma15_reg[5]  ( .D(n1854), .CK(clk), .RN(reset), .Q(sigma15[5])
         );
  DFFRHQX1 \sigma14_reg[0]  ( .D(n1836), .CK(clk), .RN(reset), .Q(sigma14[0])
         );
  DFFRHQX1 \sigma5_reg[10]  ( .D(n1768), .CK(clk), .RN(reset), .Q(sigma5[10])
         );
  DFFRHQX1 \sigma5_reg[3]  ( .D(n1761), .CK(clk), .RN(reset), .Q(sigma5[3]) );
  DFFRHQX1 \sigma7_reg[10]  ( .D(n1742), .CK(clk), .RN(reset), .Q(sigma7[10])
         );
  DFFRHQX1 \sigma1_reg[12]  ( .D(n1822), .CK(clk), .RN(reset), .Q(sigma1[12])
         );
  DFFRHQX1 \sigma15_reg[1]  ( .D(n1850), .CK(clk), .RN(reset), .Q(sigma15[1])
         );
  DFFRHQX1 \sigma8_reg[3]  ( .D(n1722), .CK(clk), .RN(reset), .Q(sigma8[3]) );
  DFFRHQX2 \sigma11_reg[7]  ( .D(n1687), .CK(clk), .RN(reset), .Q(sigma11[7])
         );
  DFFRHQX1 \sigma10_reg[0]  ( .D(n1693), .CK(clk), .RN(reset), .Q(sigma10[0])
         );
  DFFRHQX1 \sigma12_reg[5]  ( .D(n1672), .CK(clk), .RN(reset), .Q(sigma12[5])
         );
  DFFRHQX4 \sigma14_reg[6]  ( .D(n1842), .CK(clk), .RN(reset), .Q(sigma14[6])
         );
  DFFRHQX4 \sigma15_reg[8]  ( .D(n1857), .CK(clk), .RN(reset), .Q(sigma15[8])
         );
  DFFRHQX4 \sigma13_reg[4]  ( .D(n1866), .CK(clk), .RN(reset), .Q(sigma13[4])
         );
  DFFRHQX2 \sigma5_reg[0]  ( .D(n1758), .CK(clk), .RN(reset), .Q(sigma5[0]) );
  DFFRHQX4 \sigma7_reg[9]  ( .D(n1741), .CK(clk), .RN(reset), .Q(sigma7[9]) );
  DFFRHQX2 \sigma14_reg[10]  ( .D(n1846), .CK(clk), .RN(reset), .Q(sigma14[10]) );
  DFFRHQX2 \sigma1_reg[7]  ( .D(n1817), .CK(clk), .RN(reset), .Q(sigma1[7]) );
  DFFRHQX4 \sigma5_reg[11]  ( .D(n1769), .CK(clk), .RN(reset), .Q(sigma5[11])
         );
  DFFRHQX2 \sigma9_reg[1]  ( .D(n1707), .CK(clk), .RN(reset), .Q(sigma9[1]) );
  XNOR2XL U3 ( .A(L1_6[1]), .B(L1_5[1]), .Y(n433) );
  XNOR2XL U4 ( .A(L16_4[2]), .B(L16_3[2]), .Y(n543) );
  XOR2X1 U5 ( .A(n1495), .B(n1496), .Y(n1494) );
  XNOR2X1 U6 ( .A(col0[6]), .B(L5_7[6]), .Y(n1361) );
  XOR2X1 U7 ( .A(n1335), .B(n1336), .Y(n1334) );
  XNOR2X1 U8 ( .A(L9_2[10]), .B(L9_1[10]), .Y(n1336) );
  XOR2X1 U9 ( .A(n556), .B(L16_8[4]), .Y(n555) );
  XOR2X1 U10 ( .A(n557), .B(n558), .Y(n556) );
  XOR2X1 U11 ( .A(n708), .B(L14_8[10]), .Y(n707) );
  XOR2X1 U12 ( .A(n732), .B(L15_8[0]), .Y(n731) );
  XOR2X1 U13 ( .A(n796), .B(L15_8[8]), .Y(n795) );
  CLKBUFX8 U14 ( .A(col7[8]), .Y(n1904) );
  XOR2XL U15 ( .A(L13_4[11]), .B(L13_3[11]), .Y(n393) );
  XNOR2X1 U16 ( .A(L9_4[9]), .B(L9_3[9]), .Y(n871) );
  XNOR2XL U17 ( .A(L1_6[5]), .B(L1_5[5]), .Y(n465) );
  XNOR2X1 U18 ( .A(L7_2[4]), .B(L7_1[4]), .Y(n1496) );
  XNOR2X1 U19 ( .A(L7_4[4]), .B(L7_3[4]), .Y(n1495) );
  XOR2X1 U20 ( .A(n1658), .B(n1665), .Y(n678) );
  XOR2X1 U21 ( .A(L14_4[6]), .B(L14_3[6]), .Y(n1658) );
  XOR2X1 U22 ( .A(n801), .B(n802), .Y(n797) );
  XOR2X1 U23 ( .A(n1649), .B(n1650), .Y(n870) );
  XOR2X1 U24 ( .A(L13_4[4]), .B(L13_3[4]), .Y(n1649) );
  XOR2X1 U25 ( .A(n759), .B(n760), .Y(n758) );
  XNOR2X1 U26 ( .A(L15_4[3]), .B(L15_3[3]), .Y(n759) );
  XOR2X1 U27 ( .A(n1346), .B(n1361), .Y(n53) );
  XOR2X1 U28 ( .A(n490), .B(n505), .Y(n1414) );
  XOR2X1 U29 ( .A(L8_4[7]), .B(L8_3[7]), .Y(n490) );
  OAI2BB2X1 U30 ( .B0(n1331), .B1(n1914), .A0N(sigma9[10]), .A1N(n1929), .Y(
        n1716) );
  XOR2X1 U31 ( .A(n1332), .B(L9_8[10]), .Y(n1331) );
  XOR2X1 U32 ( .A(n1333), .B(n1334), .Y(n1332) );
  OAI2BB2X1 U33 ( .B0(n1491), .B1(n1916), .A0N(sigma7[4]), .A1N(n1934), .Y(
        n1736) );
  XOR2X1 U34 ( .A(n1492), .B(L7_8[4]), .Y(n1491) );
  XOR2X1 U35 ( .A(n1493), .B(n1494), .Y(n1492) );
  XOR2X1 U36 ( .A(n525), .B(n526), .Y(n524) );
  XOR2X1 U37 ( .A(n527), .B(n528), .Y(n526) );
  XOR2X1 U38 ( .A(n1893), .B(n1894), .Y(n557) );
  XOR2X1 U39 ( .A(n676), .B(L14_8[6]), .Y(n675) );
  XOR2X1 U40 ( .A(n677), .B(n678), .Y(n676) );
  XOR2X1 U41 ( .A(n709), .B(n710), .Y(n708) );
  XOR2X1 U42 ( .A(n733), .B(n734), .Y(n732) );
  XOR2X1 U43 ( .A(n797), .B(n798), .Y(n796) );
  OAI2BB2X1 U44 ( .B0(n867), .B1(n1908), .A0N(sigma13[4]), .A1N(n1940), .Y(
        n1866) );
  XOR2X1 U45 ( .A(n868), .B(L13_8[4]), .Y(n867) );
  XOR2X1 U46 ( .A(n869), .B(n870), .Y(n868) );
  CLKBUFX1 U47 ( .A(L16_1[0]), .Y(n1) );
  INVX1 U48 ( .A(sel), .Y(n9) );
  INVX1 U49 ( .A(n9), .Y(n10) );
  XNOR2XL U50 ( .A(L9_4[11]), .B(L9_3[11]), .Y(n1343) );
  XOR2X1 U51 ( .A(n524), .B(L16_8[0]), .Y(n523) );
  XNOR2XL U52 ( .A(L7_4[1]), .B(L7_3[1]), .Y(n1471) );
  XOR2XL U53 ( .A(L16_6[12]), .B(L16_5[12]), .Y(n1884) );
  XOR2XL U54 ( .A(L1_6[10]), .B(L1_5[10]), .Y(n1900) );
  XNOR2XL U55 ( .A(L1_6[11]), .B(L1_5[11]), .Y(n513) );
  INVX1 U56 ( .A(col0[1]), .Y(n17) );
  INVX1 U57 ( .A(n17), .Y(n18) );
  XNOR2XL U58 ( .A(L1_4[11]), .B(L1_3[11]), .Y(n511) );
  XNOR2XL U59 ( .A(L1_6[0]), .B(L1_5[0]), .Y(n425) );
  XNOR2X1 U60 ( .A(L2_4[11]), .B(L2_3[11]), .Y(n407) );
  INVX1 U61 ( .A(col0[6]), .Y(n20) );
  INVX1 U62 ( .A(n20), .Y(n39) );
  INVX1 U63 ( .A(col0[12]), .Y(n40) );
  INVX1 U64 ( .A(n40), .Y(n41) );
  INVX1 U65 ( .A(col0[5]), .Y(n42) );
  INVX1 U66 ( .A(n42), .Y(n47) );
  INVX1 U67 ( .A(col0[7]), .Y(n48) );
  INVX1 U68 ( .A(n48), .Y(n49) );
  INVX1 U69 ( .A(col0[9]), .Y(n50) );
  INVX1 U70 ( .A(n50), .Y(n57) );
  INVX1 U71 ( .A(col0[2]), .Y(n58) );
  INVX1 U72 ( .A(n58), .Y(n71) );
  INVX1 U73 ( .A(col0[3]), .Y(n72) );
  INVX1 U74 ( .A(n72), .Y(n129) );
  INVX1 U75 ( .A(col0[10]), .Y(n130) );
  INVX1 U76 ( .A(n130), .Y(n135) );
  INVX1 U77 ( .A(col0[11]), .Y(n136) );
  INVX1 U78 ( .A(n136), .Y(n143) );
  INVX1 U79 ( .A(col0[4]), .Y(n144) );
  INVX1 U80 ( .A(n144), .Y(n153) );
  INVX1 U81 ( .A(col0[8]), .Y(n154) );
  INVX1 U82 ( .A(n154), .Y(n161) );
  INVX1 U83 ( .A(col0[0]), .Y(n162) );
  INVX1 U84 ( .A(n162), .Y(n193) );
  XOR2XL U85 ( .A(L4_6[6]), .B(L4_5[6]), .Y(n1878) );
  XOR2X1 U86 ( .A(L13_2[4]), .B(L13_1[4]), .Y(n1650) );
  XNOR2XL U87 ( .A(L13_4[10]), .B(L13_3[10]), .Y(n919) );
  XOR2X1 U88 ( .A(L7_6[10]), .B(L7_5[10]), .Y(n1288) );
  XNOR2XL U89 ( .A(L1_4[2]), .B(L1_3[2]), .Y(n439) );
  XNOR2XL U90 ( .A(col0[3]), .B(L12_7[3]), .Y(n1215) );
  XOR2XL U91 ( .A(L12_6[3]), .B(L12_5[3]), .Y(n1208) );
  XNOR2XL U92 ( .A(L10_4[3]), .B(L10_3[3]), .Y(n1175) );
  XOR2X1 U93 ( .A(L14_4[0]), .B(L14_3[0]), .Y(n562) );
  XOR2X1 U94 ( .A(L14_2[0]), .B(L14_1[0]), .Y(n585) );
  XOR2X1 U95 ( .A(L14_4[11]), .B(L14_3[11]), .Y(n671) );
  XOR2X1 U96 ( .A(L14_2[11]), .B(L14_1[11]), .Y(n672) );
  XOR2X1 U97 ( .A(L11_4[12]), .B(L11_3[12]), .Y(n352) );
  XOR2X1 U98 ( .A(L8_4[5]), .B(L8_3[5]), .Y(n338) );
  XOR2X1 U99 ( .A(L9_4[7]), .B(L9_3[7]), .Y(n330) );
  XOR2X1 U100 ( .A(L6_4[4]), .B(L6_3[4]), .Y(n448) );
  XOR2X1 U101 ( .A(L7_4[8]), .B(L7_3[8]), .Y(n464) );
  XNOR2X1 U102 ( .A(L8_4[8]), .B(L8_3[8]), .Y(n1423) );
  XOR2X1 U103 ( .A(L8_4[9]), .B(L8_3[9]), .Y(n792) );
  XOR2X1 U104 ( .A(L4_4[4]), .B(L4_3[4]), .Y(n816) );
  XOR2X1 U105 ( .A(n1656), .B(n1657), .Y(n798) );
  XOR2X1 U106 ( .A(L15_2[8]), .B(L15_1[8]), .Y(n1657) );
  XOR2XL U107 ( .A(L6_6[4]), .B(L6_5[4]), .Y(n1896) );
  XNOR2X1 U108 ( .A(n153), .B(L6_7[4]), .Y(n1897) );
  XNOR2XL U109 ( .A(n1601), .B(L3_8[7]), .Y(n267) );
  XNOR2X1 U110 ( .A(L11_6[9]), .B(L11_5[9]), .Y(n1121) );
  XNOR2X1 U111 ( .A(L13_4[6]), .B(L13_3[6]), .Y(n887) );
  XOR2XL U112 ( .A(L15_4[11]), .B(L15_3[11]), .Y(n761) );
  XNOR2XL U113 ( .A(L5_4[7]), .B(L5_3[7]), .Y(n63) );
  XOR2XL U114 ( .A(L4_4[3]), .B(L4_3[3]), .Y(n808) );
  XNOR2XL U115 ( .A(L3_4[1]), .B(L3_3[1]), .Y(n864) );
  XOR2X1 U116 ( .A(n161), .B(L15_7[8]), .Y(n802) );
  XNOR2XL U117 ( .A(L12_4[12]), .B(L12_3[12]), .Y(n1039) );
  XOR2XL U118 ( .A(L12_4[5]), .B(L12_3[5]), .Y(n992) );
  XNOR2X1 U119 ( .A(L10_6[3]), .B(L10_5[3]), .Y(n1177) );
  XNOR2X1 U120 ( .A(L7_6[8]), .B(L7_5[8]), .Y(n1529) );
  XOR2X1 U121 ( .A(L7_6[9]), .B(L7_5[9]), .Y(n1376) );
  XOR2X1 U122 ( .A(L4_6[2]), .B(L4_5[2]), .Y(n1394) );
  XOR2X1 U123 ( .A(L12_6[4]), .B(L12_5[4]), .Y(n1402) );
  XNOR2X1 U124 ( .A(n1402), .B(n978), .Y(n973) );
  XOR2X1 U125 ( .A(L13_6[11]), .B(L13_5[11]), .Y(n1129) );
  XNOR2X1 U126 ( .A(n1129), .B(n930), .Y(n925) );
  XNOR2X1 U127 ( .A(L2_2[1]), .B(L2_1[1]), .Y(n1553) );
  XNOR2X1 U128 ( .A(n1562), .B(L12_8[11]), .Y(n1027) );
  XNOR2X1 U129 ( .A(n1592), .B(L10_8[3]), .Y(n1171) );
  XNOR2X1 U130 ( .A(n1599), .B(L13_8[7]), .Y(n891) );
  XOR2X1 U131 ( .A(n1092), .B(L11_8[6]), .Y(n1091) );
  XNOR2X1 U132 ( .A(L6_2[3]), .B(L6_1[3]), .Y(n1617) );
  XOR2X1 U133 ( .A(n559), .B(n560), .Y(n558) );
  XOR2X1 U134 ( .A(n194), .B(n217), .Y(n1206) );
  XOR2X1 U135 ( .A(L10_4[7]), .B(L10_3[7]), .Y(n194) );
  XOR2X1 U136 ( .A(L10_2[7]), .B(L10_1[7]), .Y(n217) );
  XOR2X1 U137 ( .A(n218), .B(n223), .Y(n1294) );
  XOR2X1 U138 ( .A(L9_4[5]), .B(L9_3[5]), .Y(n218) );
  XOR2X1 U139 ( .A(L9_2[5]), .B(L9_1[5]), .Y(n223) );
  XOR2X1 U140 ( .A(n224), .B(n268), .Y(n1606) );
  XOR2X1 U141 ( .A(L6_4[5]), .B(L6_3[5]), .Y(n224) );
  XOR2X1 U142 ( .A(L6_2[5]), .B(L6_1[5]), .Y(n268) );
  XOR2X1 U143 ( .A(n297), .B(n298), .Y(n1406) );
  XOR2X1 U144 ( .A(L8_4[6]), .B(L8_3[6]), .Y(n297) );
  XOR2X1 U145 ( .A(L8_2[6]), .B(L8_1[6]), .Y(n298) );
  XOR2X1 U146 ( .A(n711), .B(n712), .Y(n710) );
  XOR2X1 U147 ( .A(n327), .B(n328), .Y(n774) );
  XOR2X1 U148 ( .A(L15_4[5]), .B(L15_3[5]), .Y(n327) );
  XOR2X1 U149 ( .A(L15_2[5]), .B(L15_1[5]), .Y(n328) );
  XNOR2X1 U150 ( .A(n329), .B(n968), .Y(n966) );
  XOR2X1 U151 ( .A(L12_4[3]), .B(L12_3[3]), .Y(n329) );
  XOR2X1 U152 ( .A(n330), .B(n337), .Y(n1310) );
  XOR2X1 U153 ( .A(L9_2[7]), .B(L9_1[7]), .Y(n337) );
  XOR2X1 U154 ( .A(n338), .B(n351), .Y(n1398) );
  XOR2X1 U155 ( .A(L8_2[5]), .B(L8_1[5]), .Y(n351) );
  XNOR2XL U156 ( .A(L11_4[6]), .B(L11_3[6]), .Y(n1095) );
  XOR2X1 U157 ( .A(n352), .B(n353), .Y(n1142) );
  XOR2X1 U158 ( .A(L11_2[12]), .B(L11_1[12]), .Y(n353) );
  XOR2X1 U159 ( .A(n354), .B(n392), .Y(n1214) );
  XOR2X1 U160 ( .A(L10_4[8]), .B(L10_3[8]), .Y(n354) );
  XOR2X1 U161 ( .A(L10_2[8]), .B(L10_1[8]), .Y(n392) );
  XOR2X1 U162 ( .A(n393), .B(n394), .Y(n926) );
  XOR2X1 U163 ( .A(L13_2[11]), .B(L13_1[11]), .Y(n394) );
  XOR2X1 U164 ( .A(n396), .B(n404), .Y(n806) );
  XOR2X1 U165 ( .A(L15_4[9]), .B(L15_3[9]), .Y(n396) );
  XOR2X1 U166 ( .A(L15_2[9]), .B(L15_1[9]), .Y(n404) );
  XOR2X1 U167 ( .A(n409), .B(n410), .Y(n1374) );
  XOR2X1 U168 ( .A(L8_4[2]), .B(L8_3[2]), .Y(n409) );
  XOR2X1 U169 ( .A(L8_2[2]), .B(L8_1[2]), .Y(n410) );
  XOR2X1 U170 ( .A(n428), .B(n436), .Y(n766) );
  XOR2X1 U171 ( .A(L15_4[4]), .B(L15_3[4]), .Y(n428) );
  XOR2X1 U172 ( .A(L15_2[4]), .B(L15_1[4]), .Y(n436) );
  XOR2X1 U173 ( .A(n441), .B(n442), .Y(n670) );
  XOR2X1 U174 ( .A(L14_4[5]), .B(L14_3[5]), .Y(n441) );
  XOR2X1 U175 ( .A(L14_2[5]), .B(L14_1[5]), .Y(n442) );
  XOR2X1 U176 ( .A(n444), .B(n447), .Y(n1190) );
  XOR2X1 U177 ( .A(L10_4[5]), .B(L10_3[5]), .Y(n444) );
  XOR2X1 U178 ( .A(L10_2[5]), .B(L10_1[5]), .Y(n447) );
  XOR2X1 U179 ( .A(n448), .B(n463), .Y(n1598) );
  XOR2X1 U180 ( .A(L6_2[4]), .B(L6_1[4]), .Y(n463) );
  XOR2X1 U181 ( .A(n464), .B(n476), .Y(n1526) );
  XOR2X1 U182 ( .A(L7_2[8]), .B(L7_1[8]), .Y(n476) );
  XNOR2X1 U183 ( .A(n615), .B(n489), .Y(n614) );
  XOR2X1 U184 ( .A(L16_2[11]), .B(L16_1[11]), .Y(n489) );
  XOR2X1 U185 ( .A(L8_2[7]), .B(L8_1[7]), .Y(n505) );
  XOR2X1 U186 ( .A(n506), .B(n514), .Y(n1078) );
  XOR2X1 U187 ( .A(L11_4[4]), .B(L11_3[4]), .Y(n506) );
  XOR2X1 U188 ( .A(L11_2[4]), .B(L11_1[4]), .Y(n514) );
  XOR2X1 U189 ( .A(n516), .B(n529), .Y(n998) );
  XOR2X1 U190 ( .A(L12_4[7]), .B(L12_3[7]), .Y(n516) );
  XOR2X1 U191 ( .A(L12_2[7]), .B(L12_1[7]), .Y(n529) );
  XOR2X1 U192 ( .A(n530), .B(n545), .Y(n814) );
  XOR2X1 U193 ( .A(L15_4[10]), .B(L15_3[10]), .Y(n530) );
  XOR2X1 U194 ( .A(L15_2[10]), .B(L15_1[10]), .Y(n545) );
  XOR2X1 U195 ( .A(n546), .B(n561), .Y(n686) );
  XOR2X1 U196 ( .A(L14_4[7]), .B(L14_3[7]), .Y(n546) );
  XOR2X1 U197 ( .A(L14_2[7]), .B(L14_1[7]), .Y(n561) );
  XOR2X1 U198 ( .A(n562), .B(n585), .Y(n630) );
  XOR2X1 U199 ( .A(n586), .B(n616), .Y(n694) );
  XOR2X1 U200 ( .A(L14_4[8]), .B(L14_3[8]), .Y(n586) );
  XOR2X1 U201 ( .A(L14_2[8]), .B(L14_1[8]), .Y(n616) );
  XOR2X1 U202 ( .A(n625), .B(n626), .Y(n878) );
  XOR2X1 U203 ( .A(L13_4[5]), .B(L13_3[5]), .Y(n625) );
  XOR2X1 U204 ( .A(L13_2[5]), .B(L13_1[5]), .Y(n626) );
  XOR2X1 U205 ( .A(n631), .B(n632), .Y(n838) );
  XOR2X1 U206 ( .A(L13_4[0]), .B(L13_3[0]), .Y(n631) );
  XOR2X1 U207 ( .A(L13_2[0]), .B(L13_1[0]), .Y(n632) );
  XOR2X1 U208 ( .A(n647), .B(n648), .Y(n1102) );
  XOR2X1 U209 ( .A(L11_4[7]), .B(L11_3[7]), .Y(n647) );
  XOR2X1 U210 ( .A(L11_2[7]), .B(L11_1[7]), .Y(n648) );
  XOR2X1 U211 ( .A(n655), .B(n656), .Y(n1510) );
  XOR2X1 U212 ( .A(L7_4[6]), .B(L7_3[6]), .Y(n655) );
  XOR2X1 U213 ( .A(L7_2[6]), .B(L7_1[6]), .Y(n656) );
  XOR2X1 U214 ( .A(n663), .B(n664), .Y(n1318) );
  XOR2X1 U215 ( .A(L9_4[8]), .B(L9_3[8]), .Y(n663) );
  XOR2X1 U216 ( .A(L9_2[8]), .B(L9_1[8]), .Y(n664) );
  XOR2X1 U217 ( .A(n665), .B(n666), .Y(n990) );
  XOR2X1 U218 ( .A(L12_4[6]), .B(L12_3[6]), .Y(n665) );
  XOR2X1 U219 ( .A(L12_2[6]), .B(L12_1[6]), .Y(n666) );
  XOR2X1 U220 ( .A(n671), .B(n672), .Y(n718) );
  XOR2X1 U221 ( .A(n679), .B(n680), .Y(n902) );
  XOR2X1 U222 ( .A(L13_4[8]), .B(L13_3[8]), .Y(n679) );
  XOR2X1 U223 ( .A(L13_2[8]), .B(L13_1[8]), .Y(n680) );
  XOR2X1 U224 ( .A(n687), .B(n688), .Y(n1390) );
  XOR2X1 U225 ( .A(L8_4[4]), .B(L8_3[4]), .Y(n687) );
  XOR2X1 U226 ( .A(L8_2[4]), .B(L8_1[4]), .Y(n688) );
  XOR2X1 U227 ( .A(n695), .B(n696), .Y(n726) );
  XOR2X1 U228 ( .A(L14_4[12]), .B(L14_3[12]), .Y(n695) );
  XOR2X1 U229 ( .A(L14_2[12]), .B(L14_1[12]), .Y(n696) );
  XOR2X1 U230 ( .A(n703), .B(n704), .Y(n1086) );
  XOR2X1 U231 ( .A(L11_4[5]), .B(L11_3[5]), .Y(n703) );
  XOR2X1 U232 ( .A(L11_2[5]), .B(L11_1[5]), .Y(n704) );
  XOR2X1 U233 ( .A(n719), .B(n720), .Y(n1006) );
  XOR2X1 U234 ( .A(L12_4[8]), .B(L12_3[8]), .Y(n719) );
  XOR2X1 U235 ( .A(L12_2[8]), .B(L12_1[8]), .Y(n720) );
  XNOR2X1 U236 ( .A(n791), .B(n721), .Y(n790) );
  XOR2X1 U237 ( .A(L15_2[7]), .B(L15_1[7]), .Y(n721) );
  XOR2X1 U238 ( .A(n722), .B(n727), .Y(n1014) );
  XOR2X1 U239 ( .A(L12_4[9]), .B(L12_3[9]), .Y(n722) );
  XOR2X1 U240 ( .A(L12_2[9]), .B(L12_1[9]), .Y(n727) );
  XOR2X1 U241 ( .A(n728), .B(n736), .Y(n702) );
  XOR2X1 U242 ( .A(L14_4[9]), .B(L14_3[9]), .Y(n728) );
  XOR2X1 U243 ( .A(L14_2[9]), .B(L14_1[9]), .Y(n736) );
  XOR2X1 U244 ( .A(n761), .B(n762), .Y(n822) );
  XOR2X1 U245 ( .A(L15_2[11]), .B(L15_1[11]), .Y(n762) );
  XOR2X1 U246 ( .A(n767), .B(n768), .Y(n1046) );
  XOR2X1 U247 ( .A(L11_4[0]), .B(L11_3[0]), .Y(n767) );
  XOR2X1 U248 ( .A(L11_2[0]), .B(L11_1[0]), .Y(n768) );
  XOR2X1 U249 ( .A(n769), .B(n770), .Y(n1222) );
  XOR2X1 U250 ( .A(L10_4[9]), .B(L10_3[9]), .Y(n769) );
  XOR2X1 U251 ( .A(L10_2[9]), .B(L10_1[9]), .Y(n770) );
  XOR2X1 U252 ( .A(n775), .B(n776), .Y(n782) );
  XOR2X1 U253 ( .A(L15_4[6]), .B(L15_3[6]), .Y(n775) );
  XOR2X1 U254 ( .A(L15_2[6]), .B(L15_1[6]), .Y(n776) );
  XNOR2XL U255 ( .A(L10_4[4]), .B(L10_3[4]), .Y(n1183) );
  XOR2X1 U256 ( .A(n783), .B(n784), .Y(n1502) );
  XOR2X1 U257 ( .A(L7_4[5]), .B(L7_3[5]), .Y(n783) );
  XOR2X1 U258 ( .A(L7_2[5]), .B(L7_1[5]), .Y(n784) );
  XOR2X1 U259 ( .A(n792), .B(n799), .Y(n1430) );
  XOR2X1 U260 ( .A(L8_2[9]), .B(L8_1[9]), .Y(n799) );
  XOR2X1 U261 ( .A(n800), .B(n807), .Y(n1302) );
  XOR2X1 U262 ( .A(L9_4[6]), .B(L9_3[6]), .Y(n800) );
  XOR2X1 U263 ( .A(L9_2[6]), .B(L9_1[6]), .Y(n807) );
  XOR2X1 U264 ( .A(n808), .B(n815), .Y(n134) );
  XOR2X1 U265 ( .A(L4_2[3]), .B(L4_1[3]), .Y(n815) );
  XOR2X1 U266 ( .A(n816), .B(n823), .Y(n142) );
  XOR2X1 U267 ( .A(L4_2[4]), .B(L4_1[4]), .Y(n823) );
  XOR2X1 U268 ( .A(n824), .B(n839), .Y(n46) );
  XOR2X1 U269 ( .A(L5_4[5]), .B(L5_3[5]), .Y(n824) );
  XOR2X1 U270 ( .A(L5_2[5]), .B(L5_1[5]), .Y(n839) );
  XOR2X1 U271 ( .A(n840), .B(n847), .Y(n1518) );
  XOR2X1 U272 ( .A(L7_4[7]), .B(L7_3[7]), .Y(n840) );
  XOR2X1 U273 ( .A(L7_2[7]), .B(L7_1[7]), .Y(n847) );
  XOR2X1 U274 ( .A(n848), .B(n857), .Y(n1278) );
  XOR2X1 U275 ( .A(L9_4[3]), .B(L9_3[3]), .Y(n848) );
  XOR2X1 U276 ( .A(L9_2[3]), .B(L9_1[3]), .Y(n857) );
  XOR2X1 U277 ( .A(n858), .B(n863), .Y(n1438) );
  XOR2X1 U278 ( .A(L8_4[10]), .B(L8_3[10]), .Y(n858) );
  XOR2X1 U279 ( .A(L8_2[10]), .B(L8_1[10]), .Y(n863) );
  XOR2X1 U280 ( .A(n864), .B(n865), .Y(n222) );
  XNOR2XL U281 ( .A(L3_2[1]), .B(L3_1[1]), .Y(n865) );
  XNOR2X1 U282 ( .A(n1655), .B(n866), .Y(n38) );
  XNOR2XL U283 ( .A(L5_2[4]), .B(L5_1[4]), .Y(n866) );
  XOR2X1 U284 ( .A(n871), .B(n872), .Y(n1326) );
  XNOR2XL U285 ( .A(L9_2[9]), .B(L9_1[9]), .Y(n872) );
  XNOR2XL U286 ( .A(L1_6[3]), .B(L1_5[3]), .Y(n449) );
  XOR2X1 U287 ( .A(n879), .B(n880), .Y(n1238) );
  XOR2X1 U288 ( .A(L10_4[11]), .B(L10_3[11]), .Y(n879) );
  XOR2X1 U289 ( .A(L10_2[11]), .B(L10_1[11]), .Y(n880) );
  XNOR2X1 U290 ( .A(L9_4[10]), .B(L9_3[10]), .Y(n1335) );
  XOR2X1 U291 ( .A(L15_4[8]), .B(L15_3[8]), .Y(n1656) );
  XOR2X1 U292 ( .A(L14_2[6]), .B(L14_1[6]), .Y(n1665) );
  XNOR2X1 U293 ( .A(n735), .B(n892), .Y(n734) );
  XOR2X1 U294 ( .A(L15_2[0]), .B(L15_1[0]), .Y(n892) );
  XOR2X1 U295 ( .A(n895), .B(n896), .Y(n1557) );
  XOR2X1 U296 ( .A(L7_6[12]), .B(L7_5[12]), .Y(n895) );
  XNOR2X1 U297 ( .A(col0[12]), .B(L7_7[12]), .Y(n896) );
  XNOR2X1 U298 ( .A(n153), .B(L16_7[4]), .Y(n1894) );
  XOR2XL U299 ( .A(col0[0]), .B(L15_7[0]), .Y(n738) );
  XNOR2XL U300 ( .A(L15_6[1]), .B(L15_5[1]), .Y(n745) );
  XOR2X1 U301 ( .A(n903), .B(n904), .Y(n1365) );
  XOR2X1 U302 ( .A(L8_6[1]), .B(L8_5[1]), .Y(n903) );
  XNOR2X1 U303 ( .A(col0[1]), .B(L8_7[1]), .Y(n904) );
  XOR2X1 U304 ( .A(n913), .B(n914), .Y(n646) );
  XOR2XL U305 ( .A(L14_4[2]), .B(L14_3[2]), .Y(n913) );
  XOR2X1 U306 ( .A(L14_2[2]), .B(L14_1[2]), .Y(n914) );
  XOR2X1 U307 ( .A(n927), .B(n928), .Y(n654) );
  XOR2X1 U308 ( .A(L14_4[3]), .B(L14_3[3]), .Y(n927) );
  XOR2X1 U309 ( .A(L14_2[3]), .B(L14_1[3]), .Y(n928) );
  XOR2X1 U310 ( .A(n929), .B(n935), .Y(n1286) );
  XOR2X1 U311 ( .A(L9_4[4]), .B(L9_3[4]), .Y(n929) );
  XOR2X1 U312 ( .A(L9_2[4]), .B(L9_1[4]), .Y(n935) );
  XOR2X1 U313 ( .A(n936), .B(n945), .Y(n1478) );
  XOR2X1 U314 ( .A(L7_4[2]), .B(L7_3[2]), .Y(n936) );
  XOR2X1 U315 ( .A(L7_2[2]), .B(L7_1[2]), .Y(n945) );
  XOR2X1 U316 ( .A(n946), .B(n967), .Y(n1150) );
  XOR2X1 U317 ( .A(L10_4[0]), .B(L10_3[0]), .Y(n946) );
  XOR2X1 U318 ( .A(L10_2[0]), .B(L10_1[0]), .Y(n967) );
  XOR2X1 U319 ( .A(n969), .B(n970), .Y(n1022) );
  XOR2X1 U320 ( .A(L12_4[10]), .B(L12_3[10]), .Y(n969) );
  XOR2X1 U321 ( .A(L12_2[10]), .B(L12_1[10]), .Y(n970) );
  XOR2X1 U322 ( .A(n977), .B(n983), .Y(n934) );
  XOR2X1 U323 ( .A(L13_4[12]), .B(L13_3[12]), .Y(n977) );
  XOR2X1 U324 ( .A(L13_2[12]), .B(L13_1[12]), .Y(n983) );
  XOR2X1 U325 ( .A(n984), .B(n991), .Y(n1246) );
  XOR2X1 U326 ( .A(L10_4[12]), .B(L10_3[12]), .Y(n984) );
  XOR2X1 U327 ( .A(L10_2[12]), .B(L10_1[12]), .Y(n991) );
  XOR2X1 U328 ( .A(n992), .B(n999), .Y(n982) );
  XOR2X1 U329 ( .A(L12_2[5]), .B(L12_1[5]), .Y(n999) );
  XOR2X1 U330 ( .A(n1000), .B(n1007), .Y(n1198) );
  XOR2X1 U331 ( .A(L10_4[6]), .B(L10_3[6]), .Y(n1000) );
  XOR2X1 U332 ( .A(L10_2[6]), .B(L10_1[6]), .Y(n1007) );
  XOR2X1 U333 ( .A(n1008), .B(n1009), .Y(n1454) );
  XOR2X1 U334 ( .A(L8_4[12]), .B(L8_3[12]), .Y(n1008) );
  XOR2X1 U335 ( .A(L8_2[12]), .B(L8_1[12]), .Y(n1009) );
  XOR2X1 U336 ( .A(n1010), .B(n1015), .Y(n1270) );
  XOR2X1 U337 ( .A(L9_4[2]), .B(L9_3[2]), .Y(n1010) );
  XOR2X1 U338 ( .A(L9_2[2]), .B(L9_1[2]), .Y(n1015) );
  XOR2X1 U339 ( .A(n1016), .B(n1023), .Y(n662) );
  XOR2X1 U340 ( .A(L14_4[4]), .B(L14_3[4]), .Y(n1016) );
  XOR2X1 U341 ( .A(L14_2[4]), .B(L14_1[4]), .Y(n1023) );
  XOR2X1 U342 ( .A(n1024), .B(n1028), .Y(n1542) );
  XOR2X1 U343 ( .A(L7_4[10]), .B(L7_3[10]), .Y(n1024) );
  XOR2X1 U344 ( .A(L7_2[10]), .B(L7_1[10]), .Y(n1028) );
  XOR2X1 U345 ( .A(n1047), .B(n1048), .Y(n1070) );
  XOR2X1 U346 ( .A(L11_4[3]), .B(L11_3[3]), .Y(n1047) );
  XOR2X1 U347 ( .A(L11_2[3]), .B(L11_1[3]), .Y(n1048) );
  XOR2X1 U348 ( .A(n1049), .B(n1050), .Y(n70) );
  XOR2X1 U349 ( .A(L5_4[8]), .B(L5_3[8]), .Y(n1049) );
  XOR2X1 U350 ( .A(L5_2[8]), .B(L5_1[8]), .Y(n1050) );
  XOR2X1 U351 ( .A(L13_4[7]), .B(L13_3[7]), .Y(n1666) );
  XOR2X1 U352 ( .A(n1071), .B(n1072), .Y(n1158) );
  XOR2X1 U353 ( .A(L10_4[1]), .B(L10_3[1]), .Y(n1071) );
  XOR2X1 U354 ( .A(L10_2[1]), .B(L10_1[1]), .Y(n1072) );
  XOR2X1 U355 ( .A(n1079), .B(n1080), .Y(n1654) );
  XOR2X1 U356 ( .A(L6_4[11]), .B(L6_3[11]), .Y(n1079) );
  XOR2X1 U357 ( .A(L6_2[11]), .B(L6_1[11]), .Y(n1080) );
  XNOR2XL U358 ( .A(L3_4[2]), .B(L3_3[2]), .Y(n231) );
  XOR2X1 U359 ( .A(n1081), .B(n1082), .Y(n350) );
  XOR2X1 U360 ( .A(L2_4[4]), .B(L2_3[4]), .Y(n1081) );
  XOR2X1 U361 ( .A(L2_2[4]), .B(L2_1[4]), .Y(n1082) );
  XOR2X1 U362 ( .A(n1087), .B(n1088), .Y(n462) );
  XNOR2XL U363 ( .A(L1_4[5]), .B(L1_3[5]), .Y(n1087) );
  XNOR2X1 U364 ( .A(L1_2[5]), .B(L1_1[5]), .Y(n1088) );
  XNOR2X1 U365 ( .A(n391), .B(n1103), .Y(n390) );
  XOR2X1 U366 ( .A(L2_2[9]), .B(L2_1[9]), .Y(n1103) );
  XOR2X1 U367 ( .A(n1104), .B(n1113), .Y(n1637) );
  XOR2X1 U368 ( .A(L6_6[9]), .B(L6_5[9]), .Y(n1104) );
  XNOR2X1 U369 ( .A(n57), .B(L6_7[9]), .Y(n1113) );
  XOR2X1 U370 ( .A(n1114), .B(n1116), .Y(n13) );
  XOR2X1 U371 ( .A(L5_6[1]), .B(L5_5[1]), .Y(n1114) );
  XNOR2X1 U372 ( .A(col0[1]), .B(L5_7[1]), .Y(n1116) );
  XOR2X1 U373 ( .A(n1130), .B(n1143), .Y(n349) );
  XOR2X1 U374 ( .A(L2_6[4]), .B(L2_5[4]), .Y(n1130) );
  XNOR2X1 U375 ( .A(col0[4]), .B(L2_7[4]), .Y(n1143) );
  XOR2X1 U376 ( .A(n1144), .B(n1151), .Y(n1213) );
  XOR2X1 U377 ( .A(L10_6[8]), .B(L10_5[8]), .Y(n1144) );
  XNOR2X1 U378 ( .A(col0[8]), .B(L10_7[8]), .Y(n1151) );
  XOR2X1 U379 ( .A(n1152), .B(n1153), .Y(n1397) );
  XOR2X1 U380 ( .A(L8_6[5]), .B(L8_5[5]), .Y(n1152) );
  XNOR2X1 U381 ( .A(col0[5]), .B(L8_7[5]), .Y(n1153) );
  XOR2X1 U382 ( .A(n1154), .B(n1159), .Y(n1661) );
  XOR2X1 U383 ( .A(L6_6[12]), .B(L6_5[12]), .Y(n1154) );
  XNOR2X1 U384 ( .A(col0[12]), .B(L6_7[12]), .Y(n1159) );
  XOR2X1 U385 ( .A(n1160), .B(n1172), .Y(n5) );
  XOR2X1 U386 ( .A(L5_6[0]), .B(L5_5[0]), .Y(n1160) );
  XNOR2X1 U387 ( .A(col0[0]), .B(L5_7[0]), .Y(n1172) );
  XOR2X1 U388 ( .A(n1185), .B(n1186), .Y(n45) );
  XOR2X1 U389 ( .A(L5_6[5]), .B(L5_5[5]), .Y(n1185) );
  XNOR2X1 U390 ( .A(col0[5]), .B(L5_7[5]), .Y(n1186) );
  XOR2X1 U391 ( .A(n1191), .B(n1192), .Y(n541) );
  XOR2X1 U392 ( .A(L16_6[2]), .B(L16_5[2]), .Y(n1191) );
  XNOR2X1 U393 ( .A(col0[2]), .B(n1903), .Y(n1192) );
  XNOR2X1 U394 ( .A(n1895), .B(n1199), .Y(n765) );
  XOR2X1 U395 ( .A(n153), .B(L15_7[4]), .Y(n1199) );
  XOR2X1 U396 ( .A(n1200), .B(n1207), .Y(n1125) );
  XOR2X1 U397 ( .A(L11_6[10]), .B(L11_5[10]), .Y(n1200) );
  XNOR2X1 U398 ( .A(col0[10]), .B(L11_7[10]), .Y(n1207) );
  XOR2X1 U399 ( .A(n1208), .B(n1215), .Y(n965) );
  XOR2X1 U400 ( .A(n1216), .B(n1217), .Y(n1509) );
  XOR2X1 U401 ( .A(L7_6[6]), .B(L7_5[6]), .Y(n1216) );
  XNOR2X1 U402 ( .A(col0[6]), .B(L7_7[6]), .Y(n1217) );
  XOR2X1 U403 ( .A(n1218), .B(n1223), .Y(n861) );
  XOR2X1 U404 ( .A(L13_6[3]), .B(L13_5[3]), .Y(n1218) );
  XNOR2X1 U405 ( .A(col0[3]), .B(L13_7[3]), .Y(n1223) );
  XOR2X1 U406 ( .A(n1224), .B(n1239), .Y(n757) );
  XOR2X1 U407 ( .A(L15_6[3]), .B(L15_5[3]), .Y(n1224) );
  XNOR2X1 U408 ( .A(col0[3]), .B(L15_7[3]), .Y(n1239) );
  XOR2X1 U409 ( .A(n1240), .B(n1241), .Y(n1181) );
  XOR2X1 U410 ( .A(L10_6[4]), .B(L10_5[4]), .Y(n1240) );
  XNOR2X1 U411 ( .A(col0[4]), .B(L10_7[4]), .Y(n1241) );
  XOR2X1 U412 ( .A(n1242), .B(n1247), .Y(n853) );
  XOR2X1 U413 ( .A(L13_6[2]), .B(L13_5[2]), .Y(n1242) );
  XNOR2X1 U414 ( .A(col0[2]), .B(L13_7[2]), .Y(n1247) );
  XOR2X1 U415 ( .A(n1248), .B(n1249), .Y(n1653) );
  XOR2X1 U416 ( .A(L6_6[11]), .B(L6_5[11]), .Y(n1248) );
  XNOR2X1 U417 ( .A(col0[11]), .B(L6_7[11]), .Y(n1249) );
  XOR2X1 U418 ( .A(n1250), .B(n1265), .Y(n1429) );
  XOR2X1 U419 ( .A(L8_6[9]), .B(L8_5[9]), .Y(n1250) );
  XNOR2X1 U420 ( .A(col0[9]), .B(L8_7[9]), .Y(n1265) );
  XOR2X1 U421 ( .A(n1266), .B(n1271), .Y(n1237) );
  XOR2X1 U422 ( .A(L10_6[11]), .B(L10_5[11]), .Y(n1266) );
  XNOR2X1 U423 ( .A(col0[11]), .B(L10_7[11]), .Y(n1271) );
  XOR2XL U424 ( .A(col0[4]), .B(L3_7[4]), .Y(n250) );
  XOR2X1 U425 ( .A(n1272), .B(n1279), .Y(n1613) );
  XOR2X1 U426 ( .A(L6_6[6]), .B(L6_5[6]), .Y(n1272) );
  XNOR2X1 U427 ( .A(n39), .B(L6_7[6]), .Y(n1279) );
  XOR2X1 U428 ( .A(n1280), .B(n1287), .Y(n1549) );
  XOR2X1 U429 ( .A(L7_6[11]), .B(L7_5[11]), .Y(n1280) );
  XNOR2X1 U430 ( .A(n143), .B(L7_7[11]), .Y(n1287) );
  XOR2X1 U431 ( .A(n1288), .B(n1295), .Y(n1541) );
  XNOR2X1 U432 ( .A(col0[10]), .B(L7_7[10]), .Y(n1295) );
  XOR2X1 U433 ( .A(n1296), .B(n1303), .Y(n1461) );
  XOR2X1 U434 ( .A(L7_6[0]), .B(L7_5[0]), .Y(n1296) );
  XNOR2X1 U435 ( .A(col0[0]), .B(L7_7[0]), .Y(n1303) );
  XOR2X1 U436 ( .A(n1304), .B(n1311), .Y(n1645) );
  XOR2X1 U437 ( .A(L6_6[10]), .B(L6_5[10]), .Y(n1304) );
  XNOR2X1 U438 ( .A(n135), .B(L6_7[10]), .Y(n1311) );
  XOR2X1 U439 ( .A(n1312), .B(n1319), .Y(n1629) );
  XOR2X1 U440 ( .A(L6_6[8]), .B(L6_5[8]), .Y(n1312) );
  XNOR2X1 U441 ( .A(n161), .B(L6_7[8]), .Y(n1319) );
  XOR2X1 U442 ( .A(n1320), .B(n1327), .Y(n1605) );
  XOR2X1 U443 ( .A(L6_6[5]), .B(L6_5[5]), .Y(n1320) );
  XNOR2X1 U444 ( .A(col0[5]), .B(L6_7[5]), .Y(n1327) );
  XOR2X1 U445 ( .A(n1328), .B(n1345), .Y(n581) );
  XOR2X1 U446 ( .A(L16_6[7]), .B(L16_5[7]), .Y(n1328) );
  XNOR2X1 U447 ( .A(col0[7]), .B(L16_7[7]), .Y(n1345) );
  XOR2X1 U448 ( .A(L5_6[6]), .B(L5_5[6]), .Y(n1346) );
  XOR2X1 U449 ( .A(n1362), .B(n1369), .Y(n1517) );
  XOR2X1 U450 ( .A(L7_6[7]), .B(L7_5[7]), .Y(n1362) );
  XNOR2X1 U451 ( .A(col0[7]), .B(L7_7[7]), .Y(n1369) );
  XOR2X1 U452 ( .A(n1370), .B(n1375), .Y(n1357) );
  XOR2X1 U453 ( .A(L8_6[0]), .B(L8_5[0]), .Y(n1370) );
  XNOR2X1 U454 ( .A(n193), .B(L8_7[0]), .Y(n1375) );
  XOR2X1 U455 ( .A(n1376), .B(n1391), .Y(n1533) );
  XNOR2X1 U456 ( .A(n57), .B(L7_7[9]), .Y(n1391) );
  XOR2X1 U457 ( .A(n1392), .B(n1393), .Y(n1045) );
  XOR2X1 U458 ( .A(L11_6[0]), .B(L11_5[0]), .Y(n1392) );
  XNOR2X1 U459 ( .A(n193), .B(L11_7[0]), .Y(n1393) );
  XOR2XL U460 ( .A(col0[6]), .B(L3_7[6]), .Y(n266) );
  XOR2X1 U461 ( .A(n1394), .B(n1399), .Y(n125) );
  XNOR2X1 U462 ( .A(col0[2]), .B(L4_7[2]), .Y(n1399) );
  XOR2X1 U463 ( .A(n1400), .B(n1401), .Y(n293) );
  XOR2X1 U464 ( .A(L3_6[10]), .B(L3_5[10]), .Y(n1400) );
  XNOR2X1 U465 ( .A(col0[10]), .B(L3_7[10]), .Y(n1401) );
  XOR2X1 U466 ( .A(n1407), .B(n1408), .Y(n1389) );
  XOR2X1 U467 ( .A(L8_6[4]), .B(L8_5[4]), .Y(n1407) );
  XNOR2X1 U468 ( .A(col0[4]), .B(L8_7[4]), .Y(n1408) );
  XOR2X1 U469 ( .A(n1415), .B(n1416), .Y(n1077) );
  XOR2X1 U470 ( .A(L11_6[4]), .B(L11_5[4]), .Y(n1415) );
  XNOR2X1 U471 ( .A(n153), .B(L11_7[4]), .Y(n1416) );
  XOR2X1 U472 ( .A(n1431), .B(n1432), .Y(n189) );
  XOR2X1 U473 ( .A(L4_6[10]), .B(L4_5[10]), .Y(n1431) );
  XNOR2X1 U474 ( .A(col0[10]), .B(L4_7[10]), .Y(n1432) );
  XOR2X1 U475 ( .A(n1433), .B(n1434), .Y(n1261) );
  XOR2X1 U476 ( .A(L9_6[1]), .B(L9_5[1]), .Y(n1433) );
  XNOR2X1 U477 ( .A(n18), .B(L9_7[1]), .Y(n1434) );
  XOR2XL U478 ( .A(col0[0]), .B(L2_7[0]), .Y(n322) );
  XOR2X1 U479 ( .A(n1439), .B(n1440), .Y(n717) );
  XOR2X1 U480 ( .A(L14_6[11]), .B(L14_5[11]), .Y(n1439) );
  XNOR2XL U481 ( .A(col0[11]), .B(L14_7[11]), .Y(n1440) );
  XOR2X1 U482 ( .A(n1441), .B(n1442), .Y(n1469) );
  XOR2X1 U483 ( .A(L7_6[1]), .B(L7_5[1]), .Y(n1441) );
  XNOR2XL U484 ( .A(col0[1]), .B(L7_7[1]), .Y(n1442) );
  XOR2X1 U485 ( .A(n1455), .B(n1456), .Y(n325) );
  XOR2X1 U486 ( .A(L2_6[1]), .B(L2_5[1]), .Y(n1455) );
  XNOR2XL U487 ( .A(col0[1]), .B(L2_7[1]), .Y(n1456) );
  XOR2X1 U488 ( .A(n1465), .B(n1466), .Y(n1341) );
  XOR2X1 U489 ( .A(L9_6[11]), .B(L9_5[11]), .Y(n1465) );
  XNOR2X1 U490 ( .A(n143), .B(L9_7[11]), .Y(n1466) );
  XOR2X1 U491 ( .A(n1473), .B(n1474), .Y(n941) );
  XOR2X1 U492 ( .A(L12_6[0]), .B(L12_5[0]), .Y(n1473) );
  XNOR2XL U493 ( .A(col0[0]), .B(L12_7[0]), .Y(n1474) );
  XOR2X1 U494 ( .A(n1479), .B(n1480), .Y(n1005) );
  XOR2X1 U495 ( .A(L12_6[8]), .B(L12_5[8]), .Y(n1479) );
  XNOR2XL U496 ( .A(col0[8]), .B(L12_7[8]), .Y(n1480) );
  XOR2X1 U497 ( .A(n1489), .B(n1490), .Y(n1245) );
  XOR2X1 U498 ( .A(L10_6[12]), .B(L10_5[12]), .Y(n1489) );
  XNOR2X1 U499 ( .A(col0[12]), .B(L10_7[12]), .Y(n1490) );
  XOR2X1 U500 ( .A(n1497), .B(n1498), .Y(n1485) );
  XOR2X1 U501 ( .A(L7_6[3]), .B(L7_5[3]), .Y(n1497) );
  XNOR2XL U502 ( .A(col0[3]), .B(L7_7[3]), .Y(n1498) );
  XNOR2XL U503 ( .A(L2_6[8]), .B(L2_5[8]), .Y(n385) );
  XOR2XL U504 ( .A(col0[8]), .B(L2_7[8]), .Y(n386) );
  XOR2X1 U505 ( .A(n1503), .B(n1504), .Y(n389) );
  XOR2X1 U506 ( .A(L2_6[9]), .B(L2_5[9]), .Y(n1503) );
  XNOR2X1 U507 ( .A(col0[9]), .B(L2_7[9]), .Y(n1504) );
  XOR2X1 U508 ( .A(n1511), .B(n1512), .Y(n661) );
  XOR2X1 U509 ( .A(L14_6[4]), .B(L14_5[4]), .Y(n1511) );
  XNOR2X1 U510 ( .A(col0[4]), .B(L14_7[4]), .Y(n1512) );
  XOR2X1 U511 ( .A(n1513), .B(n1514), .Y(n1437) );
  XOR2X1 U512 ( .A(L8_6[10]), .B(L8_5[10]), .Y(n1513) );
  XNOR2XL U513 ( .A(col0[10]), .B(L8_7[10]), .Y(n1514) );
  XOR2X1 U514 ( .A(n1519), .B(n1520), .Y(n1149) );
  XNOR2X1 U515 ( .A(L10_6[0]), .B(L10_5[0]), .Y(n1519) );
  XOR2X1 U516 ( .A(n193), .B(L10_7[0]), .Y(n1520) );
  XOR2X1 U517 ( .A(n1521), .B(n1522), .Y(n1565) );
  XOR2X1 U518 ( .A(L6_6[0]), .B(L6_5[0]), .Y(n1521) );
  XNOR2X1 U519 ( .A(n193), .B(L6_7[0]), .Y(n1522) );
  XOR2X1 U520 ( .A(n1527), .B(n1528), .Y(n149) );
  XOR2X1 U521 ( .A(L4_6[5]), .B(L4_5[5]), .Y(n1527) );
  XNOR2X1 U522 ( .A(col0[5]), .B(L4_7[5]), .Y(n1528) );
  XOR2X1 U523 ( .A(n1537), .B(n1538), .Y(n485) );
  XOR2X1 U524 ( .A(L1_6[8]), .B(L1_5[8]), .Y(n1537) );
  XNOR2XL U525 ( .A(col0[8]), .B(L1_7[8]), .Y(n1538) );
  XOR2X1 U526 ( .A(n1543), .B(n1544), .Y(n525) );
  XNOR2X1 U527 ( .A(L16_6[0]), .B(L16_5[0]), .Y(n1543) );
  XOR2X1 U528 ( .A(n193), .B(L16_7[0]), .Y(n1544) );
  XNOR2X1 U529 ( .A(n1888), .B(n1545), .Y(n213) );
  XOR2X1 U530 ( .A(n193), .B(L3_7[0]), .Y(n1545) );
  XNOR2XL U531 ( .A(L2_2[2]), .B(L2_1[2]), .Y(n336) );
  XNOR2XL U532 ( .A(L1_2[10]), .B(L1_1[10]), .Y(n504) );
  XOR2X1 U533 ( .A(n1546), .B(n1553), .Y(n326) );
  XNOR2XL U534 ( .A(L2_4[1]), .B(L2_3[1]), .Y(n1546) );
  XOR2X1 U535 ( .A(n1554), .B(n1561), .Y(n446) );
  XOR2X1 U536 ( .A(L1_4[3]), .B(L1_3[3]), .Y(n1554) );
  XOR2X1 U537 ( .A(L1_2[3]), .B(L1_1[3]), .Y(n1561) );
  XNOR2XL U538 ( .A(col0[10]), .B(L1_7[10]), .Y(n1901) );
  XNOR2X1 U539 ( .A(n1029), .B(n1030), .Y(n1562) );
  XNOR2XL U540 ( .A(n1569), .B(L5_8[2]), .Y(n19) );
  XNOR2X1 U541 ( .A(n21), .B(n22), .Y(n1569) );
  XNOR2XL U542 ( .A(n1570), .B(L1_8[3]), .Y(n443) );
  XNOR2X1 U543 ( .A(n445), .B(n446), .Y(n1570) );
  XNOR2XL U544 ( .A(n1591), .B(L1_8[7]), .Y(n475) );
  XNOR2X1 U545 ( .A(n477), .B(n478), .Y(n1591) );
  XNOR2X1 U546 ( .A(n1173), .B(n1174), .Y(n1592) );
  XNOR2X1 U547 ( .A(n893), .B(n894), .Y(n1599) );
  XNOR2XL U548 ( .A(n1600), .B(L11_8[9]), .Y(n1115) );
  XNOR2X1 U549 ( .A(n1117), .B(n1118), .Y(n1600) );
  XNOR2X1 U550 ( .A(n269), .B(n270), .Y(n1601) );
  XNOR2XL U551 ( .A(n1602), .B(L2_8[10]), .Y(n395) );
  XNOR2X1 U552 ( .A(n397), .B(n398), .Y(n1602) );
  XNOR2XL U553 ( .A(n1607), .B(L2_8[11]), .Y(n403) );
  XNOR2X1 U554 ( .A(n405), .B(n406), .Y(n1607) );
  XNOR2XL U555 ( .A(n1608), .B(L1_8[1]), .Y(n427) );
  XNOR2X1 U556 ( .A(n429), .B(n430), .Y(n1608) );
  XOR2X1 U557 ( .A(n1609), .B(n1610), .Y(n862) );
  XOR2X1 U558 ( .A(L13_4[3]), .B(L13_3[3]), .Y(n1609) );
  XOR2X1 U559 ( .A(L13_2[3]), .B(L13_1[3]), .Y(n1610) );
  XNOR2X1 U560 ( .A(n1902), .B(n1617), .Y(n1590) );
  XOR2X1 U561 ( .A(n1618), .B(n1633), .Y(n909) );
  XOR2X1 U562 ( .A(L13_6[9]), .B(L13_5[9]), .Y(n1618) );
  XNOR2XL U563 ( .A(col0[9]), .B(L13_7[9]), .Y(n1633) );
  OAI2BB2X1 U564 ( .B0(n523), .B1(n1925), .A0N(sigma16[0]), .A1N(n1935), .Y(
        n1823) );
  OAI2BB2X1 U565 ( .B0(n707), .B1(n1906), .A0N(sigma14[10]), .A1N(n1937), .Y(
        n1846) );
  OAI2BB2X1 U566 ( .B0(n675), .B1(n1906), .A0N(sigma14[6]), .A1N(n1936), .Y(
        n1842) );
  OAI2BB2X1 U567 ( .B0(n795), .B1(n1908), .A0N(sigma15[8]), .A1N(n1939), .Y(
        n1857) );
  OAI2BB2X1 U568 ( .B0(n731), .B1(n1907), .A0N(sigma15[0]), .A1N(n1937), .Y(
        n1849) );
  OAI2BB2X1 U569 ( .B0(n555), .B1(n1911), .A0N(sigma16[4]), .A1N(n1929), .Y(
        n1827) );
  XNOR2XL U570 ( .A(n1634), .B(L1_8[12]), .Y(n515) );
  XNOR2X1 U571 ( .A(n517), .B(n518), .Y(n1634) );
  XNOR2XL U572 ( .A(n1641), .B(L1_8[2]), .Y(n435) );
  XNOR2X1 U573 ( .A(n437), .B(n438), .Y(n1641) );
  XNOR2X1 U574 ( .A(n513), .B(n1642), .Y(n509) );
  XNOR2XL U575 ( .A(col0[11]), .B(L1_7[11]), .Y(n1642) );
  INVX1 U576 ( .A(n1950), .Y(n1910) );
  INVX1 U577 ( .A(n1951), .Y(n1912) );
  INVX1 U578 ( .A(n1948), .Y(n1915) );
  INVX1 U579 ( .A(n1950), .Y(n1916) );
  INVX1 U580 ( .A(n1949), .Y(n1917) );
  INVX1 U581 ( .A(n1949), .Y(n1919) );
  INVX1 U582 ( .A(n1947), .Y(n1920) );
  INVX1 U583 ( .A(n1949), .Y(n1924) );
  INVX1 U584 ( .A(n1950), .Y(n1908) );
  INVX1 U585 ( .A(n1950), .Y(n1909) );
  INVX1 U586 ( .A(n1948), .Y(n1921) );
  INVX1 U587 ( .A(n1949), .Y(n1923) );
  INVX1 U588 ( .A(n1951), .Y(n1911) );
  INVX1 U589 ( .A(n1951), .Y(n1906) );
  INVX1 U590 ( .A(n1951), .Y(n1907) );
  INVX1 U591 ( .A(n1950), .Y(n1913) );
  INVX1 U593 ( .A(n1950), .Y(n1914) );
  INVX1 U594 ( .A(n1949), .Y(n1918) );
  INVX1 U595 ( .A(n1950), .Y(n1925) );
  INVX1 U596 ( .A(n1947), .Y(n1922) );
  INVX1 U597 ( .A(n1951), .Y(n1905) );
  INVX1 U598 ( .A(n1948), .Y(n1932) );
  INVX1 U599 ( .A(n1950), .Y(n1926) );
  INVX1 U600 ( .A(n1947), .Y(n1934) );
  INVX1 U601 ( .A(n1949), .Y(n1939) );
  INVX1 U602 ( .A(n1951), .Y(n1927) );
  INVX1 U603 ( .A(n1951), .Y(n1935) );
  INVX1 U604 ( .A(n1949), .Y(n1930) );
  INVX1 U605 ( .A(n1947), .Y(n1945) );
  INVX1 U606 ( .A(n1948), .Y(n1943) );
  INVX1 U607 ( .A(n1948), .Y(n1942) );
  INVX1 U608 ( .A(n1948), .Y(n1929) );
  INVX1 U609 ( .A(n1949), .Y(n1937) );
  INVX1 U610 ( .A(n1951), .Y(n1940) );
  INVX1 U611 ( .A(n1948), .Y(n1941) );
  INVX1 U612 ( .A(n1950), .Y(n1931) );
  INVX1 U613 ( .A(n1951), .Y(n1928) );
  INVX1 U614 ( .A(n1947), .Y(n1944) );
  INVX1 U615 ( .A(n1949), .Y(n1936) );
  INVX1 U616 ( .A(n1947), .Y(n1938) );
  INVX1 U617 ( .A(n1949), .Y(n1933) );
  INVX1 U618 ( .A(n1947), .Y(n1946) );
  INVX1 U619 ( .A(n3), .Y(n1951) );
  INVX1 U620 ( .A(n3), .Y(n1949) );
  INVX1 U621 ( .A(n3), .Y(n1950) );
  INVX1 U622 ( .A(n3), .Y(n1947) );
  INVX1 U623 ( .A(n3), .Y(n1948) );
  XNOR2X1 U624 ( .A(L16_2[7]), .B(L16_1[7]), .Y(n584) );
  XNOR2X1 U625 ( .A(L16_2[9]), .B(L16_1[9]), .Y(n600) );
  XNOR2X1 U626 ( .A(L16_2[12]), .B(L16_1[12]), .Y(n624) );
  XOR2X1 U627 ( .A(n1031), .B(n1032), .Y(n1030) );
  XNOR2X1 U628 ( .A(L12_2[11]), .B(L12_1[11]), .Y(n1032) );
  XNOR2X1 U629 ( .A(L12_4[11]), .B(L12_3[11]), .Y(n1031) );
  XOR2X1 U630 ( .A(n831), .B(n832), .Y(n830) );
  XNOR2X1 U631 ( .A(L15_2[12]), .B(L15_1[12]), .Y(n832) );
  XNOR2X1 U632 ( .A(L15_4[12]), .B(L15_3[12]), .Y(n831) );
  XOR2X1 U633 ( .A(n255), .B(n256), .Y(n254) );
  XNOR2X1 U634 ( .A(L3_4[5]), .B(L3_3[5]), .Y(n255) );
  XNOR2X1 U635 ( .A(L3_2[5]), .B(L3_1[5]), .Y(n256) );
  XNOR2X1 U636 ( .A(L12_6[11]), .B(L12_5[11]), .Y(n1033) );
  XNOR2XL U637 ( .A(L11_6[6]), .B(L11_5[6]), .Y(n1097) );
  XNOR2X1 U638 ( .A(L11_6[7]), .B(L11_5[7]), .Y(n1105) );
  XNOR2X1 U639 ( .A(L16_4[9]), .B(L16_3[9]), .Y(n599) );
  XNOR2X1 U640 ( .A(L16_6[11]), .B(L16_5[11]), .Y(n617) );
  XNOR2XL U641 ( .A(L12_6[12]), .B(L12_5[12]), .Y(n1041) );
  INVX1 U642 ( .A(N419), .Y(n3) );
  XOR2X1 U643 ( .A(n1343), .B(n1344), .Y(n1342) );
  XNOR2X1 U644 ( .A(L9_2[11]), .B(L9_1[11]), .Y(n1344) );
  XNOR2X1 U645 ( .A(L9_4[12]), .B(L9_3[12]), .Y(n1351) );
  XNOR2X1 U646 ( .A(L16_2[8]), .B(L16_1[8]), .Y(n592) );
  XNOR2X1 U647 ( .A(L16_2[6]), .B(L16_1[6]), .Y(n576) );
  XNOR2X1 U648 ( .A(L9_2[0]), .B(L9_1[0]), .Y(n1256) );
  XNOR2X1 U649 ( .A(L6_2[8]), .B(L6_1[8]), .Y(n1632) );
  XNOR2X1 U650 ( .A(L6_2[10]), .B(L6_1[10]), .Y(n1648) );
  XNOR2X1 U651 ( .A(L4_2[5]), .B(L4_1[5]), .Y(n152) );
  XNOR2X1 U652 ( .A(L16_2[4]), .B(L16_1[4]), .Y(n560) );
  XNOR2X1 U653 ( .A(L16_2[1]), .B(L16_1[1]), .Y(n536) );
  XNOR2X1 U654 ( .A(L16_2[2]), .B(L16_1[2]), .Y(n544) );
  XNOR2X1 U655 ( .A(L10_4[2]), .B(L10_3[2]), .Y(n1167) );
  XOR2X1 U656 ( .A(n975), .B(n976), .Y(n974) );
  XNOR2X1 U657 ( .A(L12_2[4]), .B(L12_1[4]), .Y(n976) );
  XNOR2X1 U658 ( .A(L14_2[10]), .B(L14_1[10]), .Y(n712) );
  XOR2X1 U659 ( .A(n1551), .B(n1552), .Y(n1550) );
  XNOR2X1 U660 ( .A(L7_2[11]), .B(L7_1[11]), .Y(n1552) );
  XOR2X1 U661 ( .A(n1623), .B(n1624), .Y(n1622) );
  XNOR2X1 U662 ( .A(L6_2[7]), .B(L6_1[7]), .Y(n1624) );
  XOR2X1 U663 ( .A(L5_4[4]), .B(L5_3[4]), .Y(n1655) );
  XOR2X1 U664 ( .A(n943), .B(n944), .Y(n942) );
  XNOR2X1 U665 ( .A(L12_2[0]), .B(L12_1[0]), .Y(n944) );
  XNOR2X1 U666 ( .A(L12_4[0]), .B(L12_3[0]), .Y(n943) );
  XOR2X1 U667 ( .A(n1095), .B(n1096), .Y(n1094) );
  XNOR2X1 U668 ( .A(L11_2[6]), .B(L11_1[6]), .Y(n1096) );
  XOR2X1 U669 ( .A(n1263), .B(n1264), .Y(n1262) );
  XNOR2X1 U670 ( .A(L9_2[1]), .B(L9_1[1]), .Y(n1264) );
  XNOR2X1 U671 ( .A(L9_4[1]), .B(L9_3[1]), .Y(n1263) );
  XOR2X1 U672 ( .A(n1367), .B(n1368), .Y(n1366) );
  XNOR2X1 U673 ( .A(L8_2[1]), .B(L8_1[1]), .Y(n1368) );
  XNOR2X1 U674 ( .A(L8_4[1]), .B(L8_3[1]), .Y(n1367) );
  XOR2X1 U675 ( .A(n175), .B(n176), .Y(n174) );
  XNOR2X1 U676 ( .A(L4_2[8]), .B(L4_1[8]), .Y(n176) );
  XNOR2X1 U677 ( .A(L4_4[8]), .B(L4_3[8]), .Y(n175) );
  XOR2X1 U678 ( .A(n887), .B(n888), .Y(n886) );
  XNOR2X1 U679 ( .A(L13_2[6]), .B(L13_1[6]), .Y(n888) );
  XOR2X1 U680 ( .A(n1127), .B(n1128), .Y(n1126) );
  XNOR2X1 U681 ( .A(L11_2[10]), .B(L11_1[10]), .Y(n1128) );
  XNOR2X1 U682 ( .A(L11_4[10]), .B(L11_3[10]), .Y(n1127) );
  XOR2X1 U683 ( .A(n607), .B(n608), .Y(n606) );
  XNOR2X1 U684 ( .A(L16_4[10]), .B(L16_3[10]), .Y(n607) );
  XNOR2X1 U685 ( .A(L16_2[10]), .B(L16_1[10]), .Y(n608) );
  XOR2X1 U686 ( .A(n1119), .B(n1120), .Y(n1118) );
  XNOR2X1 U687 ( .A(L11_2[9]), .B(L11_1[9]), .Y(n1120) );
  XNOR2X1 U688 ( .A(L11_4[9]), .B(L11_3[9]), .Y(n1119) );
  XOR2X1 U689 ( .A(n911), .B(n912), .Y(n910) );
  XNOR2XL U690 ( .A(L13_4[9]), .B(L13_3[9]), .Y(n911) );
  XNOR2X1 U691 ( .A(L13_2[9]), .B(L13_1[9]), .Y(n912) );
  XOR2X1 U692 ( .A(n1183), .B(n1184), .Y(n1182) );
  XNOR2X1 U693 ( .A(L10_2[4]), .B(L10_1[4]), .Y(n1184) );
  XOR2X1 U694 ( .A(n951), .B(n952), .Y(n950) );
  XNOR2X1 U695 ( .A(L12_2[1]), .B(L12_1[1]), .Y(n952) );
  XNOR2X1 U696 ( .A(L12_4[1]), .B(L12_3[1]), .Y(n951) );
  XNOR2X1 U697 ( .A(L12_2[3]), .B(L12_1[3]), .Y(n968) );
  XOR2X1 U698 ( .A(n1447), .B(n1448), .Y(n1446) );
  XNOR2X1 U699 ( .A(L8_4[11]), .B(L8_3[11]), .Y(n1447) );
  XNOR2X1 U700 ( .A(L8_2[11]), .B(L8_1[11]), .Y(n1448) );
  XOR2X1 U701 ( .A(n1639), .B(n1640), .Y(n1638) );
  XNOR2X1 U702 ( .A(L6_4[9]), .B(L6_3[9]), .Y(n1639) );
  XNOR2X1 U703 ( .A(L6_2[9]), .B(L6_1[9]), .Y(n1640) );
  XOR2X1 U704 ( .A(n79), .B(n80), .Y(n78) );
  XNOR2X1 U705 ( .A(L5_4[9]), .B(L5_3[9]), .Y(n79) );
  XNOR2X1 U706 ( .A(L5_2[9]), .B(L5_1[9]), .Y(n80) );
  XOR2X1 U707 ( .A(n367), .B(n368), .Y(n366) );
  XNOR2X1 U708 ( .A(L2_2[6]), .B(L2_1[6]), .Y(n368) );
  XNOR2X1 U709 ( .A(L2_4[6]), .B(L2_3[6]), .Y(n367) );
  XOR2X1 U710 ( .A(n855), .B(n856), .Y(n854) );
  XNOR2X1 U711 ( .A(L13_2[2]), .B(L13_1[2]), .Y(n856) );
  XNOR2X1 U712 ( .A(L13_4[2]), .B(L13_3[2]), .Y(n855) );
  XNOR2X1 U713 ( .A(L3_4[7]), .B(L3_3[7]), .Y(n271) );
  XNOR2X1 U714 ( .A(L16_4[7]), .B(L16_3[7]), .Y(n583) );
  XNOR2XL U715 ( .A(L4_4[0]), .B(L4_3[0]), .Y(n111) );
  XNOR2X1 U716 ( .A(L13_6[7]), .B(L13_5[7]), .Y(n897) );
  XNOR2X1 U717 ( .A(L6_4[12]), .B(L6_3[12]), .Y(n1663) );
  XNOR2X1 U718 ( .A(L16_4[0]), .B(L16_3[0]), .Y(n527) );
  XNOR2X1 U719 ( .A(L6_4[10]), .B(L6_3[10]), .Y(n1647) );
  XNOR2X1 U720 ( .A(L12_6[10]), .B(L12_5[10]), .Y(n1025) );
  XNOR2X1 U721 ( .A(L10_6[5]), .B(L10_5[5]), .Y(n1193) );
  XNOR2X1 U722 ( .A(L3_4[6]), .B(L3_3[6]), .Y(n263) );
  XNOR2X1 U723 ( .A(L13_6[5]), .B(L13_5[5]), .Y(n881) );
  XNOR2X1 U724 ( .A(L16_4[8]), .B(L16_3[8]), .Y(n591) );
  XNOR2X1 U725 ( .A(L16_4[12]), .B(L16_3[12]), .Y(n623) );
  XNOR2X1 U726 ( .A(L16_6[10]), .B(L16_5[10]), .Y(n609) );
  XNOR2X1 U727 ( .A(L4_4[10]), .B(L4_3[10]), .Y(n191) );
  XOR2X1 U728 ( .A(n1423), .B(n1424), .Y(n1422) );
  XNOR2X1 U729 ( .A(L8_2[8]), .B(L8_1[8]), .Y(n1424) );
  XOR2X1 U730 ( .A(n1535), .B(n1536), .Y(n1534) );
  XNOR2X1 U731 ( .A(L7_2[9]), .B(L7_1[9]), .Y(n1536) );
  XNOR2X1 U732 ( .A(L7_4[9]), .B(L7_3[9]), .Y(n1535) );
  XOR2X1 U733 ( .A(n1615), .B(n1616), .Y(n1614) );
  XNOR2X1 U734 ( .A(L6_2[6]), .B(L6_1[6]), .Y(n1616) );
  XNOR2X1 U735 ( .A(L6_4[6]), .B(L6_3[6]), .Y(n1615) );
  XOR2X1 U736 ( .A(n159), .B(n160), .Y(n158) );
  XNOR2X1 U737 ( .A(L4_2[6]), .B(L4_1[6]), .Y(n160) );
  XNOR2X1 U738 ( .A(L4_4[6]), .B(L4_3[6]), .Y(n159) );
  XNOR2X1 U739 ( .A(L7_4[0]), .B(L7_3[0]), .Y(n1463) );
  XNOR2X1 U740 ( .A(L4_4[5]), .B(L4_3[5]), .Y(n151) );
  XOR2X1 U741 ( .A(n55), .B(n56), .Y(n54) );
  XNOR2X1 U742 ( .A(L5_2[6]), .B(L5_1[6]), .Y(n56) );
  XNOR2X1 U743 ( .A(L5_4[6]), .B(L5_3[6]), .Y(n55) );
  XOR2X1 U744 ( .A(n63), .B(n64), .Y(n62) );
  XNOR2X1 U745 ( .A(L5_2[7]), .B(L5_1[7]), .Y(n64) );
  XNOR2X1 U746 ( .A(L8_4[0]), .B(L8_3[0]), .Y(n1359) );
  XNOR2X1 U747 ( .A(L4_4[1]), .B(L4_3[1]), .Y(n119) );
  XNOR2X1 U748 ( .A(L9_4[0]), .B(L9_3[0]), .Y(n1255) );
  XNOR2X1 U749 ( .A(L16_4[1]), .B(L16_3[1]), .Y(n535) );
  XNOR2X1 U750 ( .A(L16_4[5]), .B(L16_3[5]), .Y(n567) );
  XNOR2X1 U751 ( .A(L16_4[6]), .B(L16_3[6]), .Y(n575) );
  XNOR2X1 U752 ( .A(L13_6[4]), .B(L13_5[4]), .Y(n873) );
  XNOR2X1 U753 ( .A(L9_6[5]), .B(L9_5[5]), .Y(n1297) );
  XNOR2X1 U754 ( .A(L8_6[12]), .B(L8_5[12]), .Y(n1457) );
  XNOR2X1 U755 ( .A(L12_6[5]), .B(L12_5[5]), .Y(n985) );
  XNOR2X1 U756 ( .A(L11_6[5]), .B(L11_5[5]), .Y(n1089) );
  XNOR2X1 U757 ( .A(L11_6[11]), .B(L11_5[11]), .Y(n1137) );
  XNOR2X1 U758 ( .A(L13_6[10]), .B(L13_5[10]), .Y(n921) );
  XNOR2X1 U759 ( .A(L13_6[12]), .B(L13_5[12]), .Y(n937) );
  XNOR2X1 U760 ( .A(L11_6[12]), .B(L11_5[12]), .Y(n1145) );
  XNOR2X1 U761 ( .A(L9_6[4]), .B(L9_5[4]), .Y(n1289) );
  XOR2X1 U762 ( .A(n1135), .B(n1136), .Y(n1134) );
  XNOR2X1 U763 ( .A(L11_2[11]), .B(L11_1[11]), .Y(n1136) );
  XNOR2X1 U764 ( .A(L11_4[11]), .B(L11_3[11]), .Y(n1135) );
  XNOR2X1 U765 ( .A(L5_2[1]), .B(L5_1[1]), .Y(n16) );
  XNOR2XL U766 ( .A(L5_4[1]), .B(L5_3[1]), .Y(n15) );
  XNOR2X1 U767 ( .A(L3_2[7]), .B(L3_1[7]), .Y(n272) );
  XNOR2X1 U768 ( .A(L4_2[1]), .B(L4_1[1]), .Y(n120) );
  XNOR2X1 U769 ( .A(L6_2[2]), .B(L6_1[2]), .Y(n1584) );
  XNOR2X1 U770 ( .A(L2_4[2]), .B(L2_3[2]), .Y(n335) );
  XOR2X1 U771 ( .A(n745), .B(n746), .Y(n741) );
  XOR2X1 U772 ( .A(n18), .B(L15_7[1]), .Y(n746) );
  XOR2X1 U773 ( .A(n369), .B(n370), .Y(n365) );
  XNOR2X1 U774 ( .A(L2_6[6]), .B(L2_5[6]), .Y(n369) );
  XOR2X1 U775 ( .A(n777), .B(n778), .Y(n773) );
  XNOR2X1 U776 ( .A(L15_6[5]), .B(L15_5[5]), .Y(n777) );
  XOR2X1 U777 ( .A(n87), .B(n88), .Y(n86) );
  XNOR2X1 U778 ( .A(L5_2[10]), .B(L5_1[10]), .Y(n88) );
  XOR2X1 U779 ( .A(n793), .B(n794), .Y(n789) );
  XOR2X1 U780 ( .A(L15_7[7]), .B(col0[7]), .Y(n794) );
  XOR2X1 U781 ( .A(n95), .B(n96), .Y(n94) );
  XNOR2X1 U782 ( .A(L5_2[11]), .B(L5_1[11]), .Y(n96) );
  XOR2X1 U783 ( .A(n577), .B(n578), .Y(n573) );
  XNOR2X1 U784 ( .A(L16_6[6]), .B(L16_5[6]), .Y(n577) );
  XOR2X1 U785 ( .A(n39), .B(L16_7[6]), .Y(n578) );
  XNOR2X1 U786 ( .A(L6_2[0]), .B(L6_1[0]), .Y(n1568) );
  XOR2X1 U787 ( .A(n135), .B(L12_7[10]), .Y(n1026) );
  XOR2X1 U788 ( .A(n753), .B(n754), .Y(n749) );
  XOR2X1 U789 ( .A(n71), .B(L15_7[2]), .Y(n754) );
  XOR2X1 U790 ( .A(n71), .B(L8_7[2]), .Y(n1378) );
  XNOR2X1 U791 ( .A(L9_2[12]), .B(L9_1[12]), .Y(n1352) );
  XNOR2X1 U792 ( .A(L8_2[0]), .B(L8_1[0]), .Y(n1360) );
  XNOR2X1 U793 ( .A(L7_2[0]), .B(L7_1[0]), .Y(n1464) );
  XNOR2X1 U794 ( .A(L7_2[12]), .B(L7_1[12]), .Y(n1560) );
  XNOR2X1 U795 ( .A(L6_2[12]), .B(L6_1[12]), .Y(n1664) );
  XNOR2X1 U796 ( .A(L5_2[12]), .B(L5_1[12]), .Y(n104) );
  XNOR2X1 U797 ( .A(L4_2[10]), .B(L4_1[10]), .Y(n192) );
  XNOR2X1 U798 ( .A(L10_2[2]), .B(L10_1[2]), .Y(n1168) );
  XNOR2X1 U799 ( .A(L6_2[1]), .B(L6_1[1]), .Y(n1576) );
  XOR2X1 U800 ( .A(n639), .B(n640), .Y(n638) );
  XNOR2X1 U801 ( .A(L14_4[1]), .B(L14_3[1]), .Y(n639) );
  XNOR2X1 U802 ( .A(L14_2[1]), .B(L14_1[1]), .Y(n640) );
  XNOR2X1 U803 ( .A(L16_2[5]), .B(L16_1[5]), .Y(n568) );
  XOR2X1 U804 ( .A(n135), .B(L13_7[10]), .Y(n922) );
  XOR2X1 U805 ( .A(n431), .B(n432), .Y(n430) );
  XNOR2X1 U806 ( .A(L1_2[1]), .B(L1_1[1]), .Y(n432) );
  XOR2X1 U807 ( .A(n167), .B(n168), .Y(n166) );
  XNOR2X1 U808 ( .A(L4_2[7]), .B(L4_1[7]), .Y(n168) );
  XOR2X1 U809 ( .A(n47), .B(L10_7[5]), .Y(n1194) );
  XOR2X1 U810 ( .A(n247), .B(n248), .Y(n246) );
  XNOR2X1 U811 ( .A(L3_2[4]), .B(L3_1[4]), .Y(n248) );
  XOR2X1 U812 ( .A(n1063), .B(n1064), .Y(n1062) );
  XNOR2X1 U813 ( .A(L11_2[2]), .B(L11_1[2]), .Y(n1064) );
  XOR2X1 U814 ( .A(n1666), .B(n1875), .Y(n894) );
  XOR2X1 U815 ( .A(L13_2[7]), .B(L13_1[7]), .Y(n1875) );
  XOR2X1 U816 ( .A(n1876), .B(n1877), .Y(n846) );
  XOR2XL U817 ( .A(L13_4[1]), .B(L13_3[1]), .Y(n1876) );
  XOR2X1 U818 ( .A(L13_2[1]), .B(L13_1[1]), .Y(n1877) );
  XOR2X1 U819 ( .A(n71), .B(L7_7[2]), .Y(n1482) );
  XOR2X1 U820 ( .A(n135), .B(L16_7[10]), .Y(n610) );
  XOR2X1 U821 ( .A(n129), .B(L16_7[3]), .Y(n554) );
  XOR2X1 U822 ( .A(n49), .B(L8_7[7]), .Y(n1418) );
  XOR2X1 U823 ( .A(n1878), .B(n1879), .Y(n157) );
  XNOR2X1 U824 ( .A(col0[6]), .B(L4_7[6]), .Y(n1879) );
  XOR2X1 U825 ( .A(n249), .B(n250), .Y(n245) );
  XNOR2X1 U826 ( .A(L3_6[4]), .B(L3_5[4]), .Y(n249) );
  XOR2X1 U827 ( .A(n41), .B(L12_7[12]), .Y(n1042) );
  XOR2X1 U828 ( .A(n143), .B(L11_7[11]), .Y(n1138) );
  XOR2X1 U829 ( .A(col0[4]), .B(L9_7[4]), .Y(n1290) );
  XOR2X1 U830 ( .A(col0[9]), .B(L11_7[9]), .Y(n1122) );
  XOR2X1 U831 ( .A(n49), .B(L11_7[7]), .Y(n1106) );
  XOR2X1 U832 ( .A(n41), .B(L8_7[12]), .Y(n1458) );
  XOR2X1 U833 ( .A(n41), .B(L15_7[12]), .Y(n834) );
  XOR2X1 U834 ( .A(n265), .B(n266), .Y(n261) );
  XNOR2X1 U835 ( .A(L3_6[6]), .B(L3_5[6]), .Y(n265) );
  XOR2X1 U836 ( .A(n71), .B(L11_7[2]), .Y(n1066) );
  XOR2X1 U837 ( .A(n1039), .B(n1040), .Y(n1038) );
  XNOR2X1 U838 ( .A(L12_2[12]), .B(L12_1[12]), .Y(n1040) );
  XOR2X1 U839 ( .A(n1073), .B(n1074), .Y(n1069) );
  XNOR2X1 U840 ( .A(L11_6[3]), .B(L11_5[3]), .Y(n1073) );
  XOR2X1 U841 ( .A(n129), .B(L11_7[3]), .Y(n1074) );
  XOR2X1 U842 ( .A(n1111), .B(n1112), .Y(n1110) );
  XNOR2X1 U843 ( .A(L11_2[8]), .B(L11_1[8]), .Y(n1112) );
  XNOR2X1 U844 ( .A(L11_4[8]), .B(L11_3[8]), .Y(n1111) );
  XOR2X1 U845 ( .A(n1383), .B(n1384), .Y(n1382) );
  XNOR2X1 U846 ( .A(L8_2[3]), .B(L8_1[3]), .Y(n1384) );
  XNOR2X1 U847 ( .A(L8_4[3]), .B(L8_3[3]), .Y(n1383) );
  XOR2X1 U848 ( .A(n751), .B(n752), .Y(n750) );
  XNOR2X1 U849 ( .A(L15_2[2]), .B(L15_1[2]), .Y(n752) );
  XNOR2X1 U850 ( .A(L15_4[2]), .B(L15_3[2]), .Y(n751) );
  XOR2X1 U851 ( .A(n919), .B(n920), .Y(n918) );
  XNOR2X1 U852 ( .A(L13_2[10]), .B(L13_1[10]), .Y(n920) );
  XOR2X1 U853 ( .A(n1487), .B(n1488), .Y(n1486) );
  XNOR2X1 U854 ( .A(L7_4[3]), .B(L7_3[3]), .Y(n1487) );
  XNOR2X1 U855 ( .A(L7_2[3]), .B(L7_1[3]), .Y(n1488) );
  XOR2X1 U856 ( .A(n7), .B(n8), .Y(n6) );
  XNOR2X1 U857 ( .A(L5_2[0]), .B(L5_1[0]), .Y(n8) );
  XNOR2X1 U858 ( .A(L5_4[0]), .B(L5_3[0]), .Y(n7) );
  XOR2X1 U859 ( .A(n127), .B(n128), .Y(n126) );
  XNOR2X1 U860 ( .A(L4_2[2]), .B(L4_1[2]), .Y(n128) );
  XNOR2X1 U861 ( .A(L4_4[2]), .B(L4_3[2]), .Y(n127) );
  XOR2X1 U862 ( .A(n183), .B(n184), .Y(n182) );
  XNOR2X1 U863 ( .A(L4_2[9]), .B(L4_1[9]), .Y(n184) );
  XNOR2X1 U864 ( .A(L4_4[9]), .B(L4_3[9]), .Y(n183) );
  XOR2X1 U865 ( .A(n199), .B(n200), .Y(n198) );
  XNOR2X1 U866 ( .A(L4_2[11]), .B(L4_1[11]), .Y(n200) );
  XNOR2X1 U867 ( .A(L4_4[11]), .B(L4_3[11]), .Y(n199) );
  XOR2X1 U868 ( .A(n231), .B(n232), .Y(n230) );
  XNOR2X1 U869 ( .A(L3_2[2]), .B(L3_1[2]), .Y(n232) );
  XOR2X1 U870 ( .A(n279), .B(n280), .Y(n278) );
  XNOR2X1 U871 ( .A(L3_2[8]), .B(L3_1[8]), .Y(n280) );
  XNOR2X1 U872 ( .A(L3_4[8]), .B(L3_3[8]), .Y(n279) );
  XOR2X1 U873 ( .A(n303), .B(n304), .Y(n302) );
  XNOR2X1 U874 ( .A(L3_2[11]), .B(L3_1[11]), .Y(n304) );
  XNOR2X1 U875 ( .A(L3_4[11]), .B(L3_3[11]), .Y(n303) );
  XOR2X1 U876 ( .A(n359), .B(n360), .Y(n358) );
  XNOR2X1 U877 ( .A(L2_4[5]), .B(L2_3[5]), .Y(n359) );
  XNOR2X1 U878 ( .A(L2_2[5]), .B(L2_1[5]), .Y(n360) );
  XOR2X1 U879 ( .A(n375), .B(n376), .Y(n374) );
  XNOR2X1 U880 ( .A(L2_2[7]), .B(L2_1[7]), .Y(n376) );
  XNOR2X1 U881 ( .A(L2_4[7]), .B(L2_3[7]), .Y(n375) );
  XOR2X1 U882 ( .A(n383), .B(n384), .Y(n382) );
  XNOR2X1 U883 ( .A(L2_2[8]), .B(L2_1[8]), .Y(n384) );
  XNOR2X1 U884 ( .A(L2_4[8]), .B(L2_3[8]), .Y(n383) );
  XOR2X1 U885 ( .A(n455), .B(n456), .Y(n454) );
  XNOR2X1 U886 ( .A(L1_2[4]), .B(L1_1[4]), .Y(n456) );
  XNOR2X1 U887 ( .A(L1_4[4]), .B(L1_3[4]), .Y(n455) );
  XOR2X1 U888 ( .A(n551), .B(n552), .Y(n550) );
  XNOR2XL U889 ( .A(L16_4[3]), .B(L16_3[3]), .Y(n551) );
  XNOR2X1 U890 ( .A(L16_2[3]), .B(L16_1[3]), .Y(n552) );
  XOR2X1 U891 ( .A(n743), .B(n744), .Y(n742) );
  XNOR2X1 U892 ( .A(L15_2[1]), .B(L15_1[1]), .Y(n744) );
  XNOR2X1 U893 ( .A(L15_4[1]), .B(L15_3[1]), .Y(n743) );
  XNOR2X1 U894 ( .A(L8_6[2]), .B(L8_5[2]), .Y(n1377) );
  XOR2X1 U895 ( .A(n41), .B(L11_7[12]), .Y(n1146) );
  XOR2X1 U896 ( .A(n143), .B(L16_7[11]), .Y(n618) );
  XOR2X1 U897 ( .A(n143), .B(L12_7[11]), .Y(n1034) );
  XOR2X1 U898 ( .A(col0[6]), .B(L11_7[6]), .Y(n1098) );
  XOR2X1 U899 ( .A(col0[5]), .B(L9_7[5]), .Y(n1298) );
  XOR2X1 U900 ( .A(n153), .B(L13_7[4]), .Y(n874) );
  XOR2X1 U901 ( .A(n473), .B(n474), .Y(n469) );
  XNOR2X1 U902 ( .A(L1_6[6]), .B(L1_5[6]), .Y(n473) );
  XOR2X1 U903 ( .A(n39), .B(L1_7[6]), .Y(n474) );
  XNOR2X1 U904 ( .A(L12_4[2]), .B(L12_3[2]), .Y(n959) );
  XNOR2X1 U905 ( .A(L15_6[12]), .B(L15_5[12]), .Y(n833) );
  XNOR2X1 U906 ( .A(L15_6[0]), .B(L15_5[0]), .Y(n737) );
  XNOR2X1 U907 ( .A(L3_4[12]), .B(L3_3[12]), .Y(n311) );
  XOR2X1 U908 ( .A(n295), .B(n296), .Y(n294) );
  XNOR2X1 U909 ( .A(L3_2[10]), .B(L3_1[10]), .Y(n296) );
  XNOR2X1 U910 ( .A(L3_4[10]), .B(L3_3[10]), .Y(n295) );
  XNOR2X1 U911 ( .A(L8_6[7]), .B(L8_5[7]), .Y(n1417) );
  XNOR2X1 U912 ( .A(L4_4[12]), .B(L4_3[12]), .Y(n207) );
  XOR2X1 U913 ( .A(n287), .B(n288), .Y(n286) );
  XNOR2X1 U914 ( .A(L3_2[9]), .B(L3_1[9]), .Y(n288) );
  XNOR2X1 U915 ( .A(L3_4[9]), .B(L3_3[9]), .Y(n287) );
  XNOR2X1 U916 ( .A(L6_4[2]), .B(L6_3[2]), .Y(n1583) );
  XNOR2X1 U917 ( .A(L5_4[12]), .B(L5_3[12]), .Y(n103) );
  XOR2X1 U918 ( .A(n1161), .B(n1162), .Y(n1157) );
  XOR2X1 U919 ( .A(n18), .B(L10_7[1]), .Y(n1162) );
  XNOR2X1 U920 ( .A(L10_6[1]), .B(L10_5[1]), .Y(n1161) );
  XOR2X1 U921 ( .A(n25), .B(n26), .Y(n21) );
  XOR2X1 U922 ( .A(col0[2]), .B(L5_7[2]), .Y(n26) );
  XNOR2X1 U923 ( .A(L5_6[2]), .B(L5_5[2]), .Y(n25) );
  XNOR2X1 U924 ( .A(L13_6[8]), .B(L13_5[8]), .Y(n905) );
  XOR2X1 U925 ( .A(n1471), .B(n1472), .Y(n1470) );
  XNOR2X1 U926 ( .A(L7_2[1]), .B(L7_1[1]), .Y(n1472) );
  XOR2X1 U927 ( .A(n233), .B(n234), .Y(n229) );
  XOR2X1 U928 ( .A(n71), .B(L3_7[2]), .Y(n234) );
  XNOR2X1 U929 ( .A(L3_6[2]), .B(L3_5[2]), .Y(n233) );
  XOR2X1 U930 ( .A(n641), .B(n642), .Y(n637) );
  XOR2X1 U931 ( .A(n18), .B(L14_7[1]), .Y(n642) );
  XNOR2XL U932 ( .A(L14_6[1]), .B(L14_5[1]), .Y(n641) );
  XNOR2XL U933 ( .A(L6_4[1]), .B(L6_3[1]), .Y(n1575) );
  XOR2X1 U934 ( .A(n1055), .B(n1056), .Y(n1054) );
  XNOR2X1 U935 ( .A(L11_2[1]), .B(L11_1[1]), .Y(n1056) );
  XNOR2X1 U936 ( .A(L11_4[1]), .B(L11_3[1]), .Y(n1055) );
  XNOR2X1 U937 ( .A(L11_6[2]), .B(L11_5[2]), .Y(n1065) );
  XNOR2X1 U938 ( .A(L16_4[4]), .B(L16_3[4]), .Y(n559) );
  XOR2X1 U939 ( .A(n1880), .B(n1881), .Y(n1493) );
  XOR2X1 U940 ( .A(L7_6[4]), .B(L7_5[4]), .Y(n1880) );
  XNOR2XL U941 ( .A(col0[4]), .B(L7_7[4]), .Y(n1881) );
  XOR2X1 U942 ( .A(n1505), .B(n1506), .Y(n1501) );
  XOR2X1 U943 ( .A(col0[5]), .B(L7_7[5]), .Y(n1506) );
  XNOR2X1 U944 ( .A(L7_6[5]), .B(L7_5[5]), .Y(n1505) );
  XOR2X1 U945 ( .A(n257), .B(n258), .Y(n253) );
  XOR2X1 U946 ( .A(n47), .B(L3_7[5]), .Y(n258) );
  XNOR2X1 U947 ( .A(L3_6[5]), .B(L3_5[5]), .Y(n257) );
  XOR2X1 U948 ( .A(n313), .B(n314), .Y(n309) );
  XOR2X1 U949 ( .A(n41), .B(L3_7[12]), .Y(n314) );
  XNOR2X1 U950 ( .A(L3_6[12]), .B(L3_5[12]), .Y(n313) );
  XOR2X1 U951 ( .A(n1882), .B(n1883), .Y(n37) );
  XOR2X1 U952 ( .A(L5_6[4]), .B(L5_5[4]), .Y(n1882) );
  XNOR2X1 U953 ( .A(n153), .B(L5_7[4]), .Y(n1883) );
  XNOR2X1 U954 ( .A(L7_6[2]), .B(L7_5[2]), .Y(n1481) );
  XOR2X1 U955 ( .A(n1231), .B(n1232), .Y(n1230) );
  XNOR2X1 U956 ( .A(L10_2[10]), .B(L10_1[10]), .Y(n1232) );
  XNOR2X1 U957 ( .A(L10_4[10]), .B(L10_3[10]), .Y(n1231) );
  XOR2X1 U958 ( .A(n649), .B(n650), .Y(n645) );
  XOR2X1 U959 ( .A(n71), .B(L14_7[2]), .Y(n650) );
  XOR2X1 U960 ( .A(n97), .B(n98), .Y(n93) );
  XOR2X1 U961 ( .A(n143), .B(L5_7[11]), .Y(n98) );
  XOR2X1 U962 ( .A(n1884), .B(n1885), .Y(n621) );
  XNOR2XL U963 ( .A(col0[12]), .B(L16_7[12]), .Y(n1885) );
  XOR2X1 U964 ( .A(n1886), .B(n1887), .Y(n405) );
  XOR2X1 U965 ( .A(L2_6[11]), .B(L2_5[11]), .Y(n1886) );
  XNOR2X1 U966 ( .A(col0[11]), .B(L2_7[11]), .Y(n1887) );
  XOR2X1 U967 ( .A(n465), .B(n466), .Y(n461) );
  XNOR2X1 U968 ( .A(L12_2[2]), .B(L12_1[2]), .Y(n960) );
  XOR2X1 U969 ( .A(n31), .B(n32), .Y(n30) );
  XNOR2X1 U970 ( .A(L5_2[3]), .B(L5_1[3]), .Y(n32) );
  XNOR2XL U971 ( .A(L5_4[3]), .B(L5_3[3]), .Y(n31) );
  XOR2X1 U972 ( .A(n239), .B(n240), .Y(n238) );
  XNOR2XL U973 ( .A(L3_2[3]), .B(L3_1[3]), .Y(n240) );
  XNOR2XL U974 ( .A(L3_4[3]), .B(L3_3[3]), .Y(n239) );
  XOR2X1 U975 ( .A(n105), .B(n106), .Y(n101) );
  XNOR2X1 U976 ( .A(L5_6[12]), .B(L5_5[12]), .Y(n105) );
  XOR2X1 U977 ( .A(n41), .B(L5_7[12]), .Y(n106) );
  XOR2X1 U978 ( .A(n601), .B(n602), .Y(n597) );
  XNOR2X1 U979 ( .A(L16_6[9]), .B(L16_5[9]), .Y(n601) );
  XOR2X1 U980 ( .A(col0[9]), .B(L16_7[9]), .Y(n602) );
  XOR2X1 U981 ( .A(n1585), .B(n1586), .Y(n1581) );
  XNOR2X1 U982 ( .A(L6_6[2]), .B(L6_5[2]), .Y(n1585) );
  XOR2X1 U983 ( .A(L3_6[0]), .B(L3_5[0]), .Y(n1888) );
  XOR2X1 U984 ( .A(n785), .B(n786), .Y(n781) );
  XNOR2X1 U985 ( .A(L15_6[6]), .B(L15_5[6]), .Y(n785) );
  XOR2X1 U986 ( .A(n1889), .B(n1890), .Y(n1109) );
  XOR2X1 U987 ( .A(L11_6[8]), .B(L11_5[8]), .Y(n1889) );
  XNOR2XL U988 ( .A(col0[8]), .B(L11_7[8]), .Y(n1890) );
  XOR2X1 U989 ( .A(n729), .B(n730), .Y(n725) );
  XNOR2X1 U990 ( .A(L14_6[12]), .B(L14_5[12]), .Y(n729) );
  XOR2X1 U991 ( .A(n1449), .B(n1450), .Y(n1445) );
  XNOR2X1 U992 ( .A(L8_6[11]), .B(L8_5[11]), .Y(n1449) );
  XOR2X1 U993 ( .A(n1891), .B(n1892), .Y(n333) );
  XOR2X1 U994 ( .A(L2_6[2]), .B(L2_5[2]), .Y(n1891) );
  XNOR2XL U995 ( .A(col0[2]), .B(L2_7[2]), .Y(n1892) );
  XOR2X1 U996 ( .A(n417), .B(n418), .Y(n413) );
  XNOR2X1 U997 ( .A(L2_6[12]), .B(L2_5[12]), .Y(n417) );
  XOR2X1 U998 ( .A(n1001), .B(n1002), .Y(n997) );
  XOR2X1 U999 ( .A(n49), .B(L12_7[7]), .Y(n1002) );
  XNOR2X1 U1000 ( .A(L12_6[7]), .B(L12_5[7]), .Y(n1001) );
  XOR2X1 U1001 ( .A(n1337), .B(n1338), .Y(n1333) );
  XNOR2X1 U1002 ( .A(L9_6[10]), .B(L9_5[10]), .Y(n1337) );
  XOR2X1 U1003 ( .A(n135), .B(L9_7[10]), .Y(n1338) );
  XOR2X1 U1004 ( .A(L16_6[4]), .B(L16_5[4]), .Y(n1893) );
  XOR2X1 U1005 ( .A(n953), .B(n954), .Y(n949) );
  XNOR2X1 U1006 ( .A(L12_6[1]), .B(L12_5[1]), .Y(n953) );
  XOR2X1 U1007 ( .A(n18), .B(L12_7[1]), .Y(n954) );
  XOR2X1 U1008 ( .A(n1057), .B(n1058), .Y(n1053) );
  XOR2X1 U1009 ( .A(n18), .B(L11_7[1]), .Y(n1058) );
  XNOR2X1 U1010 ( .A(L11_6[1]), .B(L11_5[1]), .Y(n1057) );
  XOR2X1 U1011 ( .A(n1177), .B(n1178), .Y(n1173) );
  XOR2X1 U1012 ( .A(col0[3]), .B(L10_7[3]), .Y(n1178) );
  XOR2X1 U1013 ( .A(n1209), .B(n1210), .Y(n1205) );
  XNOR2X1 U1014 ( .A(L10_6[7]), .B(L10_5[7]), .Y(n1209) );
  XOR2X1 U1015 ( .A(n49), .B(L10_7[7]), .Y(n1210) );
  XOR2X1 U1016 ( .A(n1257), .B(n1258), .Y(n1253) );
  XNOR2X1 U1017 ( .A(L9_6[0]), .B(L9_5[0]), .Y(n1257) );
  XOR2X1 U1018 ( .A(n193), .B(L9_7[0]), .Y(n1258) );
  XOR2X1 U1019 ( .A(n1273), .B(n1274), .Y(n1269) );
  XNOR2X1 U1020 ( .A(L9_6[2]), .B(L9_5[2]), .Y(n1273) );
  XOR2X1 U1021 ( .A(col0[2]), .B(L9_7[2]), .Y(n1274) );
  XOR2X1 U1022 ( .A(n1529), .B(n1530), .Y(n1525) );
  XOR2X1 U1023 ( .A(n161), .B(L7_7[8]), .Y(n1530) );
  XOR2X1 U1024 ( .A(n1577), .B(n1578), .Y(n1573) );
  XOR2XL U1025 ( .A(col0[1]), .B(L6_7[1]), .Y(n1578) );
  XNOR2X1 U1026 ( .A(L6_6[1]), .B(L6_5[1]), .Y(n1577) );
  XOR2X1 U1027 ( .A(n1593), .B(n1594), .Y(n1589) );
  XNOR2X1 U1028 ( .A(L6_6[3]), .B(L6_5[3]), .Y(n1593) );
  XOR2X1 U1029 ( .A(n129), .B(L6_7[3]), .Y(n1594) );
  XOR2X1 U1030 ( .A(n113), .B(n114), .Y(n109) );
  XNOR2X1 U1031 ( .A(L4_6[0]), .B(L4_5[0]), .Y(n113) );
  XOR2X1 U1032 ( .A(n193), .B(L4_7[0]), .Y(n114) );
  XOR2X1 U1033 ( .A(n121), .B(n122), .Y(n117) );
  XOR2X1 U1034 ( .A(col0[1]), .B(L4_7[1]), .Y(n122) );
  XNOR2X1 U1035 ( .A(L4_6[1]), .B(L4_5[1]), .Y(n121) );
  XOR2X1 U1036 ( .A(n177), .B(n178), .Y(n173) );
  XNOR2X1 U1037 ( .A(L4_6[8]), .B(L4_5[8]), .Y(n177) );
  XOR2X1 U1038 ( .A(n161), .B(L4_7[8]), .Y(n178) );
  XOR2X1 U1039 ( .A(n201), .B(n202), .Y(n197) );
  XNOR2X1 U1040 ( .A(L4_6[11]), .B(L4_5[11]), .Y(n201) );
  XOR2X1 U1041 ( .A(n143), .B(L4_7[11]), .Y(n202) );
  XOR2X1 U1042 ( .A(n209), .B(n210), .Y(n205) );
  XOR2X1 U1043 ( .A(n41), .B(L4_7[12]), .Y(n210) );
  XNOR2X1 U1044 ( .A(L4_6[12]), .B(L4_5[12]), .Y(n209) );
  XOR2X1 U1045 ( .A(n305), .B(n306), .Y(n301) );
  XNOR2X1 U1046 ( .A(L3_6[11]), .B(L3_5[11]), .Y(n305) );
  XOR2X1 U1047 ( .A(n143), .B(L3_7[11]), .Y(n306) );
  XOR2X1 U1048 ( .A(n377), .B(n378), .Y(n373) );
  XNOR2X1 U1049 ( .A(L2_6[7]), .B(L2_5[7]), .Y(n377) );
  XOR2X1 U1050 ( .A(n49), .B(L2_7[7]), .Y(n378) );
  XOR2X1 U1051 ( .A(n537), .B(n538), .Y(n533) );
  XNOR2X1 U1052 ( .A(L16_6[1]), .B(L16_5[1]), .Y(n537) );
  XOR2X1 U1053 ( .A(n18), .B(L16_7[1]), .Y(n538) );
  XOR2X1 U1054 ( .A(n569), .B(n570), .Y(n565) );
  XNOR2X1 U1055 ( .A(L16_6[5]), .B(L16_5[5]), .Y(n569) );
  XOR2X1 U1056 ( .A(n47), .B(L16_7[5]), .Y(n570) );
  XOR2X1 U1057 ( .A(n593), .B(n594), .Y(n589) );
  XNOR2X1 U1058 ( .A(L16_6[8]), .B(L16_5[8]), .Y(n593) );
  XOR2X1 U1059 ( .A(n161), .B(L16_7[8]), .Y(n594) );
  XOR2X1 U1060 ( .A(n633), .B(n634), .Y(n629) );
  XOR2X1 U1061 ( .A(n193), .B(L14_7[0]), .Y(n634) );
  XNOR2X1 U1062 ( .A(L14_6[0]), .B(L14_5[0]), .Y(n633) );
  XOR2X1 U1063 ( .A(L15_6[4]), .B(L15_5[4]), .Y(n1895) );
  XOR2X1 U1064 ( .A(n809), .B(n810), .Y(n805) );
  XNOR2X1 U1065 ( .A(L15_6[9]), .B(L15_5[9]), .Y(n809) );
  XOR2X1 U1066 ( .A(col0[9]), .B(L15_7[9]), .Y(n810) );
  XOR2X1 U1067 ( .A(n1625), .B(n1626), .Y(n1621) );
  XOR2X1 U1068 ( .A(n49), .B(L6_7[7]), .Y(n1626) );
  XNOR2X1 U1069 ( .A(L6_6[7]), .B(L6_5[7]), .Y(n1625) );
  XOR2X1 U1070 ( .A(n1353), .B(n1354), .Y(n1349) );
  XOR2X1 U1071 ( .A(n41), .B(L9_7[12]), .Y(n1354) );
  XNOR2X1 U1072 ( .A(L9_6[12]), .B(L9_5[12]), .Y(n1353) );
  XOR2X1 U1073 ( .A(n1409), .B(n1410), .Y(n1405) );
  XNOR2X1 U1074 ( .A(L8_6[6]), .B(L8_5[6]), .Y(n1409) );
  XOR2X1 U1075 ( .A(n39), .B(L8_7[6]), .Y(n1410) );
  XOR2X1 U1076 ( .A(n1896), .B(n1897), .Y(n1597) );
  XOR2X1 U1077 ( .A(n1305), .B(n1306), .Y(n1301) );
  XNOR2X1 U1078 ( .A(L9_6[6]), .B(L9_5[6]), .Y(n1305) );
  XOR2X1 U1079 ( .A(col0[6]), .B(L9_7[6]), .Y(n1306) );
  XOR2X1 U1080 ( .A(n1201), .B(n1202), .Y(n1197) );
  XNOR2X1 U1081 ( .A(L10_6[6]), .B(L10_5[6]), .Y(n1201) );
  XOR2X1 U1082 ( .A(n39), .B(L10_7[6]), .Y(n1202) );
  XOR2X1 U1083 ( .A(n65), .B(n66), .Y(n61) );
  XOR2X1 U1084 ( .A(n49), .B(L5_7[7]), .Y(n66) );
  XNOR2X1 U1085 ( .A(L5_6[7]), .B(L5_5[7]), .Y(n65) );
  XOR2X1 U1086 ( .A(n1321), .B(n1322), .Y(n1317) );
  XOR2X1 U1087 ( .A(col0[8]), .B(L9_7[8]), .Y(n1322) );
  XNOR2X1 U1088 ( .A(L9_6[8]), .B(L9_5[8]), .Y(n1321) );
  XOR2X1 U1089 ( .A(n145), .B(n146), .Y(n141) );
  XOR2X1 U1090 ( .A(L4_7[4]), .B(n153), .Y(n146) );
  XNOR2X1 U1091 ( .A(L4_6[4]), .B(L4_5[4]), .Y(n145) );
  XOR2X1 U1092 ( .A(n1385), .B(n1386), .Y(n1381) );
  XOR2X1 U1093 ( .A(n129), .B(L8_7[3]), .Y(n1386) );
  XNOR2X1 U1094 ( .A(L8_6[3]), .B(L8_5[3]), .Y(n1385) );
  XOR2X1 U1095 ( .A(n169), .B(n170), .Y(n165) );
  XNOR2X1 U1096 ( .A(L4_6[7]), .B(L4_5[7]), .Y(n169) );
  XOR2X1 U1097 ( .A(n49), .B(L4_7[7]), .Y(n170) );
  XOR2X1 U1098 ( .A(n74), .B(n73), .Y(n69) );
  XNOR2X1 U1099 ( .A(L5_6[8]), .B(L5_5[8]), .Y(n73) );
  XOR2X1 U1100 ( .A(n161), .B(L5_7[8]), .Y(n74) );
  XOR2X1 U1101 ( .A(n657), .B(n658), .Y(n653) );
  XNOR2X1 U1102 ( .A(L14_6[3]), .B(L14_5[3]), .Y(n657) );
  XOR2X1 U1103 ( .A(n129), .B(L14_7[3]), .Y(n658) );
  XOR2X1 U1104 ( .A(n81), .B(n82), .Y(n77) );
  XNOR2X1 U1105 ( .A(L5_6[9]), .B(L5_5[9]), .Y(n81) );
  XOR2X1 U1106 ( .A(n57), .B(L5_7[9]), .Y(n82) );
  XOR2X1 U1107 ( .A(n993), .B(n994), .Y(n989) );
  XOR2X1 U1108 ( .A(n39), .B(L12_7[6]), .Y(n994) );
  XNOR2X1 U1109 ( .A(L12_6[6]), .B(L12_5[6]), .Y(n993) );
  XOR2X1 U1110 ( .A(n89), .B(n90), .Y(n85) );
  XOR2X1 U1111 ( .A(n135), .B(L5_7[10]), .Y(n90) );
  XNOR2X1 U1112 ( .A(L5_6[10]), .B(L5_5[10]), .Y(n89) );
  XOR2X1 U1113 ( .A(n961), .B(n962), .Y(n957) );
  XOR2X1 U1114 ( .A(n71), .B(L12_7[2]), .Y(n962) );
  XNOR2X1 U1115 ( .A(L12_6[2]), .B(L12_5[2]), .Y(n961) );
  XOR2X1 U1116 ( .A(n1017), .B(n1018), .Y(n1013) );
  XOR2X1 U1117 ( .A(n57), .B(L12_7[9]), .Y(n1018) );
  XNOR2X1 U1118 ( .A(L12_6[9]), .B(L12_5[9]), .Y(n1017) );
  XOR2X1 U1119 ( .A(n1169), .B(n1170), .Y(n1165) );
  XOR2X1 U1120 ( .A(n71), .B(L10_7[2]), .Y(n1170) );
  XNOR2X1 U1121 ( .A(L10_6[2]), .B(L10_5[2]), .Y(n1169) );
  XOR2X1 U1122 ( .A(n1225), .B(n1226), .Y(n1221) );
  XNOR2X1 U1123 ( .A(L10_6[9]), .B(L10_5[9]), .Y(n1225) );
  XOR2X1 U1124 ( .A(n57), .B(L10_7[9]), .Y(n1226) );
  XOR2X1 U1125 ( .A(n1233), .B(n1234), .Y(n1229) );
  XOR2X1 U1126 ( .A(n135), .B(L10_7[10]), .Y(n1234) );
  XNOR2X1 U1127 ( .A(L10_6[10]), .B(L10_5[10]), .Y(n1233) );
  XOR2X1 U1128 ( .A(n1281), .B(n1282), .Y(n1277) );
  XOR2X1 U1129 ( .A(col0[3]), .B(L9_7[3]), .Y(n1282) );
  XNOR2X1 U1130 ( .A(L9_6[3]), .B(L9_5[3]), .Y(n1281) );
  XOR2X1 U1131 ( .A(n1313), .B(n1314), .Y(n1309) );
  XOR2X1 U1132 ( .A(col0[7]), .B(L9_7[7]), .Y(n1314) );
  XNOR2X1 U1133 ( .A(L9_6[7]), .B(L9_5[7]), .Y(n1313) );
  XOR2X1 U1134 ( .A(n1425), .B(n1426), .Y(n1421) );
  XNOR2X1 U1135 ( .A(L8_6[8]), .B(L8_5[8]), .Y(n1425) );
  XOR2X1 U1136 ( .A(n161), .B(L8_7[8]), .Y(n1426) );
  XOR2X1 U1137 ( .A(n33), .B(n34), .Y(n29) );
  XOR2X1 U1138 ( .A(n129), .B(L5_7[3]), .Y(n34) );
  XNOR2X1 U1139 ( .A(L5_6[3]), .B(L5_5[3]), .Y(n33) );
  XOR2X1 U1140 ( .A(n137), .B(n138), .Y(n133) );
  XOR2X1 U1141 ( .A(n129), .B(L4_7[3]), .Y(n138) );
  XNOR2X1 U1142 ( .A(L4_6[3]), .B(L4_5[3]), .Y(n137) );
  XOR2X1 U1143 ( .A(n185), .B(n186), .Y(n181) );
  XNOR2X1 U1144 ( .A(L4_6[9]), .B(L4_5[9]), .Y(n185) );
  XOR2X1 U1145 ( .A(n57), .B(L4_7[9]), .Y(n186) );
  XOR2X1 U1146 ( .A(n225), .B(n226), .Y(n221) );
  XNOR2X1 U1147 ( .A(L3_6[1]), .B(L3_5[1]), .Y(n225) );
  XOR2X1 U1148 ( .A(n18), .B(L3_7[1]), .Y(n226) );
  XOR2X1 U1149 ( .A(n241), .B(n242), .Y(n237) );
  XOR2X1 U1150 ( .A(n129), .B(L3_7[3]), .Y(n242) );
  XNOR2XL U1151 ( .A(L3_6[3]), .B(L3_5[3]), .Y(n241) );
  XOR2X1 U1152 ( .A(n273), .B(n274), .Y(n269) );
  XOR2X1 U1153 ( .A(col0[7]), .B(L3_7[7]), .Y(n274) );
  XNOR2X1 U1154 ( .A(L3_6[7]), .B(L3_5[7]), .Y(n273) );
  XOR2X1 U1155 ( .A(n281), .B(n282), .Y(n277) );
  XNOR2X1 U1156 ( .A(L3_6[8]), .B(L3_5[8]), .Y(n281) );
  XOR2X1 U1157 ( .A(n161), .B(L3_7[8]), .Y(n282) );
  XOR2X1 U1158 ( .A(n289), .B(n290), .Y(n285) );
  XOR2X1 U1159 ( .A(n57), .B(L3_7[9]), .Y(n290) );
  XNOR2X1 U1160 ( .A(L3_6[9]), .B(L3_5[9]), .Y(n289) );
  XOR2X1 U1161 ( .A(n321), .B(n322), .Y(n317) );
  XNOR2X1 U1162 ( .A(L2_6[0]), .B(L2_5[0]), .Y(n321) );
  XOR2X1 U1163 ( .A(n345), .B(n346), .Y(n341) );
  XOR2X1 U1164 ( .A(n129), .B(L2_7[3]), .Y(n346) );
  XNOR2X1 U1165 ( .A(L2_6[3]), .B(L2_5[3]), .Y(n345) );
  XOR2X1 U1166 ( .A(n361), .B(n362), .Y(n357) );
  XNOR2X1 U1167 ( .A(L2_6[5]), .B(L2_5[5]), .Y(n361) );
  XOR2X1 U1168 ( .A(n47), .B(L2_7[5]), .Y(n362) );
  XOR2X1 U1169 ( .A(n385), .B(n386), .Y(n381) );
  XOR2X1 U1170 ( .A(n401), .B(n402), .Y(n397) );
  XOR2XL U1171 ( .A(col0[10]), .B(L2_7[10]), .Y(n402) );
  XNOR2X1 U1172 ( .A(L2_6[10]), .B(L2_5[10]), .Y(n401) );
  XOR2X1 U1173 ( .A(n457), .B(n458), .Y(n453) );
  XNOR2X1 U1174 ( .A(L1_6[4]), .B(L1_5[4]), .Y(n457) );
  XOR2X1 U1175 ( .A(n153), .B(L1_7[4]), .Y(n458) );
  XOR2X1 U1176 ( .A(n481), .B(n482), .Y(n477) );
  XOR2X1 U1177 ( .A(col0[7]), .B(L1_7[7]), .Y(n482) );
  XNOR2X1 U1178 ( .A(L1_6[7]), .B(L1_5[7]), .Y(n481) );
  XOR2X1 U1179 ( .A(n673), .B(n674), .Y(n669) );
  XNOR2X1 U1180 ( .A(L14_6[5]), .B(L14_5[5]), .Y(n673) );
  XOR2X1 U1181 ( .A(n47), .B(L14_7[5]), .Y(n674) );
  XOR2X1 U1182 ( .A(n681), .B(n682), .Y(n677) );
  XNOR2X1 U1183 ( .A(L14_6[6]), .B(L14_5[6]), .Y(n681) );
  XOR2X1 U1184 ( .A(n39), .B(L14_7[6]), .Y(n682) );
  XOR2X1 U1185 ( .A(n689), .B(n690), .Y(n685) );
  XNOR2X1 U1186 ( .A(L14_6[7]), .B(L14_5[7]), .Y(n689) );
  XOR2X1 U1187 ( .A(n49), .B(L14_7[7]), .Y(n690) );
  XOR2X1 U1188 ( .A(n697), .B(n698), .Y(n693) );
  XOR2X1 U1189 ( .A(n161), .B(L14_7[8]), .Y(n698) );
  XNOR2X1 U1190 ( .A(L14_6[8]), .B(L14_5[8]), .Y(n697) );
  XOR2X1 U1191 ( .A(n705), .B(n706), .Y(n701) );
  XOR2X1 U1192 ( .A(col0[9]), .B(L14_7[9]), .Y(n706) );
  XNOR2X1 U1193 ( .A(L14_6[9]), .B(L14_5[9]), .Y(n705) );
  XOR2X1 U1194 ( .A(n713), .B(n714), .Y(n709) );
  XOR2X1 U1195 ( .A(n135), .B(L14_7[10]), .Y(n714) );
  XNOR2X1 U1196 ( .A(L14_6[10]), .B(L14_5[10]), .Y(n713) );
  XOR2X1 U1197 ( .A(n817), .B(n818), .Y(n813) );
  XNOR2X1 U1198 ( .A(L15_6[10]), .B(L15_5[10]), .Y(n817) );
  XOR2X1 U1199 ( .A(n135), .B(L15_7[10]), .Y(n818) );
  XOR2X1 U1200 ( .A(n825), .B(n826), .Y(n821) );
  XOR2X1 U1201 ( .A(n143), .B(L15_7[11]), .Y(n826) );
  XNOR2X1 U1202 ( .A(L15_6[11]), .B(L15_5[11]), .Y(n825) );
  XOR2X1 U1203 ( .A(n841), .B(n842), .Y(n837) );
  XOR2XL U1204 ( .A(col0[0]), .B(L13_7[0]), .Y(n842) );
  XNOR2X1 U1205 ( .A(L13_6[0]), .B(L13_5[0]), .Y(n841) );
  XOR2X1 U1206 ( .A(n849), .B(n850), .Y(n845) );
  XOR2X1 U1207 ( .A(n18), .B(L13_7[1]), .Y(n850) );
  XNOR2XL U1208 ( .A(L13_6[1]), .B(L13_5[1]), .Y(n849) );
  XOR2X1 U1209 ( .A(n889), .B(n890), .Y(n885) );
  XOR2X1 U1210 ( .A(n39), .B(L13_7[6]), .Y(n890) );
  XNOR2X1 U1211 ( .A(L13_6[6]), .B(L13_5[6]), .Y(n889) );
  XOR2X1 U1212 ( .A(n1329), .B(n1330), .Y(n1325) );
  XOR2X1 U1213 ( .A(n57), .B(L9_7[9]), .Y(n1330) );
  XNOR2X1 U1214 ( .A(L9_6[9]), .B(L9_5[9]), .Y(n1329) );
  XNOR2X1 U1215 ( .A(L3_2[6]), .B(L3_1[6]), .Y(n264) );
  XOR2X1 U1216 ( .A(n47), .B(L11_7[5]), .Y(n1090) );
  XOR2X1 U1217 ( .A(n1898), .B(n1899), .Y(n437) );
  XOR2X1 U1218 ( .A(L1_6[2]), .B(L1_5[2]), .Y(n1898) );
  XNOR2XL U1219 ( .A(col0[2]), .B(L1_7[2]), .Y(n1899) );
  XNOR2X1 U1220 ( .A(L4_2[0]), .B(L4_1[0]), .Y(n112) );
  XNOR2X1 U1221 ( .A(L3_2[12]), .B(L3_1[12]), .Y(n312) );
  XNOR2X1 U1222 ( .A(L2_2[11]), .B(L2_1[11]), .Y(n408) );
  XOR2X1 U1223 ( .A(n503), .B(n504), .Y(n502) );
  XNOR2X1 U1224 ( .A(L1_4[10]), .B(L1_3[10]), .Y(n503) );
  XNOR2X1 U1225 ( .A(L5_2[2]), .B(L5_1[2]), .Y(n24) );
  XNOR2X1 U1226 ( .A(L1_2[6]), .B(L4_1[12]), .Y(n208) );
  XNOR2X1 U1227 ( .A(L2_2[10]), .B(L2_1[10]), .Y(n400) );
  XOR2X1 U1228 ( .A(n495), .B(n496), .Y(n494) );
  XNOR2X1 U1229 ( .A(L1_2[9]), .B(L2_1[10]), .Y(n496) );
  XOR2X1 U1230 ( .A(col0[1]), .B(L1_7[1]), .Y(n434) );
  XOR2X1 U1231 ( .A(col0[7]), .B(L13_7[7]), .Y(n898) );
  XOR2XL U1232 ( .A(col0[8]), .B(L13_7[8]), .Y(n906) );
  XOR2X1 U1233 ( .A(n343), .B(n344), .Y(n342) );
  XNOR2X1 U1234 ( .A(L2_2[3]), .B(L2_1[3]), .Y(n344) );
  XNOR2XL U1235 ( .A(L2_4[3]), .B(L2_3[3]), .Y(n343) );
  XOR2X1 U1236 ( .A(n471), .B(n472), .Y(n470) );
  XNOR2X1 U1237 ( .A(L1_2[6]), .B(L1_1[6]), .Y(n472) );
  XNOR2X1 U1238 ( .A(L1_4[6]), .B(L1_3[6]), .Y(n471) );
  XOR2X1 U1239 ( .A(n487), .B(n488), .Y(n486) );
  XNOR2X1 U1240 ( .A(L1_4[8]), .B(L1_3[8]), .Y(n487) );
  XNOR2X1 U1241 ( .A(L1_2[8]), .B(L1_1[8]), .Y(n488) );
  XNOR2X1 U1242 ( .A(L2_4[10]), .B(L2_3[10]), .Y(n399) );
  XNOR2X1 U1243 ( .A(L1_4[7]), .B(L1_3[7]), .Y(n479) );
  XOR2X1 U1244 ( .A(n1900), .B(n1901), .Y(n501) );
  XNOR2X1 U1245 ( .A(L1_2[7]), .B(L1_1[7]), .Y(n480) );
  XOR2XL U1246 ( .A(col0[0]), .B(L1_7[0]), .Y(n426) );
  XOR2X1 U1247 ( .A(n117), .B(n118), .Y(n116) );
  XOR2X1 U1248 ( .A(n119), .B(n120), .Y(n118) );
  XOR2X1 U1249 ( .A(n596), .B(L16_8[9]), .Y(n595) );
  XOR2X1 U1250 ( .A(n597), .B(n598), .Y(n596) );
  XOR2X1 U1251 ( .A(n599), .B(n600), .Y(n598) );
  XOR2X1 U1252 ( .A(n572), .B(L16_8[6]), .Y(n571) );
  XOR2X1 U1253 ( .A(n573), .B(n574), .Y(n572) );
  XOR2X1 U1254 ( .A(n575), .B(n576), .Y(n574) );
  XOR2X1 U1255 ( .A(n433), .B(n434), .Y(n429) );
  XOR2X1 U1256 ( .A(n1285), .B(n1286), .Y(n1284) );
  XOR2X1 U1257 ( .A(n1289), .B(n1290), .Y(n1285) );
  XOR2X1 U1258 ( .A(n1245), .B(n1246), .Y(n1244) );
  OAI2BB2X1 U1259 ( .B0(n539), .B1(n1925), .A0N(sigma16[2]), .A1N(n1935), .Y(
        n1825) );
  XOR2X1 U1260 ( .A(n540), .B(L16_8[2]), .Y(n539) );
  XOR2X1 U1261 ( .A(n541), .B(n542), .Y(n540) );
  XOR2X1 U1262 ( .A(n543), .B(n544), .Y(n542) );
  OAI2BB2X1 U1263 ( .B0(n611), .B1(n1905), .A0N(sigma16[11]), .A1N(n1935), .Y(
        n1834) );
  XOR2X1 U1264 ( .A(n612), .B(L16_8[11]), .Y(n611) );
  XOR2X1 U1265 ( .A(n613), .B(n614), .Y(n612) );
  XOR2X1 U1266 ( .A(n617), .B(n618), .Y(n613) );
  OAI2BB2X1 U1267 ( .B0(n1067), .B1(n1911), .A0N(sigma11[3]), .A1N(n1944), .Y(
        n1683) );
  XOR2X1 U1268 ( .A(n1068), .B(L11_8[3]), .Y(n1067) );
  XOR2X1 U1269 ( .A(n1069), .B(n1070), .Y(n1068) );
  OAI2BB2X1 U1270 ( .B0(n91), .B1(n1923), .A0N(sigma5[11]), .A1N(n1933), .Y(
        n1769) );
  XOR2X1 U1271 ( .A(n92), .B(L5_8[11]), .Y(n91) );
  XOR2X1 U1272 ( .A(n93), .B(n94), .Y(n92) );
  OAI2BB2X1 U1273 ( .B0(n787), .B1(n1907), .A0N(sigma15[7]), .A1N(n1938), .Y(
        n1856) );
  XOR2X1 U1274 ( .A(n788), .B(L15_8[7]), .Y(n787) );
  XOR2X1 U1275 ( .A(n789), .B(n790), .Y(n788) );
  OAI2BB2X1 U1276 ( .B0(n1627), .B1(n1918), .A0N(sigma6[8]), .A1N(n1928), .Y(
        n1753) );
  XOR2X1 U1277 ( .A(n1628), .B(L6_8[8]), .Y(n1627) );
  XOR2X1 U1278 ( .A(n1629), .B(n1630), .Y(n1628) );
  XOR2X1 U1279 ( .A(n1631), .B(n1632), .Y(n1630) );
  OAI2BB2X1 U1280 ( .B0(n651), .B1(n1906), .A0N(sigma14[3]), .A1N(n1936), .Y(
        n1839) );
  XOR2X1 U1281 ( .A(n652), .B(L14_8[3]), .Y(n651) );
  XOR2X1 U1282 ( .A(n653), .B(n654), .Y(n652) );
  OAI2BB2X1 U1283 ( .B0(n363), .B1(n1921), .A0N(sigma2[6]), .A1N(n1941), .Y(
        n1803) );
  XOR2X1 U1284 ( .A(n364), .B(L2_8[6]), .Y(n363) );
  XOR2X1 U1285 ( .A(n365), .B(n366), .Y(n364) );
  OAI2BB2X1 U1286 ( .B0(n947), .B1(n1909), .A0N(sigma12[1]), .A1N(n1942), .Y(
        n1668) );
  XOR2X1 U1287 ( .A(n948), .B(L12_8[1]), .Y(n947) );
  XOR2X1 U1288 ( .A(n949), .B(n950), .Y(n948) );
  OAI2BB2X1 U1289 ( .B0(n963), .B1(n1910), .A0N(sigma12[3]), .A1N(n1942), .Y(
        n1670) );
  XOR2X1 U1290 ( .A(n964), .B(L12_8[3]), .Y(n963) );
  XOR2X1 U1291 ( .A(n965), .B(n966), .Y(n964) );
  OAI2BB2X1 U1292 ( .B0(n1027), .B1(n1910), .A0N(sigma12[11]), .A1N(n1943), 
        .Y(n1678) );
  XOR2X1 U1293 ( .A(n1033), .B(n1034), .Y(n1029) );
  OAI2BB2X1 U1294 ( .B0(n1035), .B1(n1911), .A0N(sigma12[12]), .A1N(n1943), 
        .Y(n1679) );
  XOR2X1 U1295 ( .A(n1036), .B(L12_8[12]), .Y(n1035) );
  XOR2X1 U1296 ( .A(n1037), .B(n1038), .Y(n1036) );
  XOR2X1 U1297 ( .A(n1041), .B(n1042), .Y(n1037) );
  OAI2BB2X1 U1298 ( .B0(n1051), .B1(n1911), .A0N(sigma11[1]), .A1N(n1943), .Y(
        n1681) );
  XOR2X1 U1299 ( .A(n1052), .B(L11_8[1]), .Y(n1051) );
  XOR2X1 U1300 ( .A(n1053), .B(n1054), .Y(n1052) );
  OAI2BB2X1 U1301 ( .B0(n1059), .B1(n1911), .A0N(sigma11[2]), .A1N(n1944), .Y(
        n1682) );
  XOR2X1 U1302 ( .A(n1060), .B(L11_8[2]), .Y(n1059) );
  XOR2X1 U1303 ( .A(n1061), .B(n1062), .Y(n1060) );
  XOR2X1 U1304 ( .A(n1065), .B(n1066), .Y(n1061) );
  OAI2BB2X1 U1305 ( .B0(n1091), .B1(n1911), .A0N(sigma11[6]), .A1N(n1944), .Y(
        n1686) );
  XOR2X1 U1306 ( .A(n1093), .B(n1094), .Y(n1092) );
  XOR2X1 U1307 ( .A(n1097), .B(n1098), .Y(n1093) );
  OAI2BB2X1 U1308 ( .B0(n1107), .B1(n1912), .A0N(sigma11[8]), .A1N(n1945), .Y(
        n1688) );
  XOR2X1 U1309 ( .A(n1108), .B(L11_8[8]), .Y(n1107) );
  XOR2X1 U1310 ( .A(n1109), .B(n1110), .Y(n1108) );
  OAI2BB2X1 U1311 ( .B0(n1155), .B1(n1912), .A0N(sigma10[1]), .A1N(n1945), .Y(
        n1694) );
  XOR2X1 U1312 ( .A(n1156), .B(L10_8[1]), .Y(n1155) );
  XOR2X1 U1313 ( .A(n1157), .B(n1158), .Y(n1156) );
  OAI2BB2X1 U1314 ( .B0(n1171), .B1(n1912), .A0N(sigma10[3]), .A1N(n1946), .Y(
        n1696) );
  XOR2X1 U1315 ( .A(n1175), .B(n1176), .Y(n1174) );
  OAI2BB2X1 U1316 ( .B0(n1187), .B1(n1913), .A0N(sigma10[5]), .A1N(n1946), .Y(
        n1698) );
  XOR2X1 U1317 ( .A(n1188), .B(L10_8[5]), .Y(n1187) );
  XOR2X1 U1318 ( .A(n1189), .B(n1190), .Y(n1188) );
  XOR2X1 U1319 ( .A(n1193), .B(n1194), .Y(n1189) );
  OAI2BB2X1 U1320 ( .B0(n1203), .B1(n1913), .A0N(sigma10[7]), .A1N(n1927), .Y(
        n1700) );
  XOR2X1 U1321 ( .A(n1204), .B(L10_8[7]), .Y(n1203) );
  XOR2X1 U1322 ( .A(n1205), .B(n1206), .Y(n1204) );
  OAI2BB2X1 U1323 ( .B0(n1211), .B1(n1913), .A0N(sigma10[8]), .A1N(n1926), .Y(
        n1701) );
  XOR2X1 U1324 ( .A(n1212), .B(L10_8[8]), .Y(n1211) );
  XOR2X1 U1325 ( .A(n1213), .B(n1214), .Y(n1212) );
  OAI2BB2X1 U1326 ( .B0(n1259), .B1(n1913), .A0N(sigma9[1]), .A1N(n1926), .Y(
        n1707) );
  XOR2X1 U1327 ( .A(n1260), .B(L9_8[1]), .Y(n1259) );
  XOR2X1 U1328 ( .A(n1261), .B(n1262), .Y(n1260) );
  OAI2BB2X1 U1329 ( .B0(n1307), .B1(n1914), .A0N(sigma9[7]), .A1N(n1928), .Y(
        n1713) );
  XOR2X1 U1330 ( .A(n1308), .B(L9_8[7]), .Y(n1307) );
  XOR2X1 U1331 ( .A(n1309), .B(n1310), .Y(n1308) );
  OAI2BB2X1 U1332 ( .B0(n1323), .B1(n1914), .A0N(sigma9[9]), .A1N(n1929), .Y(
        n1715) );
  XOR2X1 U1333 ( .A(n1324), .B(L9_8[9]), .Y(n1323) );
  XOR2X1 U1334 ( .A(n1325), .B(n1326), .Y(n1324) );
  OAI2BB2X1 U1335 ( .B0(n1363), .B1(n1915), .A0N(sigma8[1]), .A1N(n1930), .Y(
        n1720) );
  XOR2X1 U1336 ( .A(n1364), .B(L8_8[1]), .Y(n1363) );
  XOR2X1 U1337 ( .A(n1365), .B(n1366), .Y(n1364) );
  OAI2BB2X1 U1338 ( .B0(n1371), .B1(n1915), .A0N(sigma8[2]), .A1N(n1930), .Y(
        n1721) );
  XOR2X1 U1339 ( .A(n1372), .B(L8_8[2]), .Y(n1371) );
  XOR2X1 U1340 ( .A(n1373), .B(n1374), .Y(n1372) );
  XOR2X1 U1341 ( .A(n1377), .B(n1378), .Y(n1373) );
  OAI2BB2X1 U1342 ( .B0(n1435), .B1(n1916), .A0N(sigma8[10]), .A1N(n1932), .Y(
        n1729) );
  XOR2X1 U1343 ( .A(n1436), .B(L8_8[10]), .Y(n1435) );
  XOR2X1 U1344 ( .A(n1437), .B(n1438), .Y(n1436) );
  OAI2BB2X1 U1345 ( .B0(n1475), .B1(n1916), .A0N(sigma7[2]), .A1N(n1933), .Y(
        n1734) );
  XOR2X1 U1346 ( .A(n1476), .B(L7_8[2]), .Y(n1475) );
  XOR2X1 U1347 ( .A(n1477), .B(n1478), .Y(n1476) );
  XOR2X1 U1348 ( .A(n1481), .B(n1482), .Y(n1477) );
  OAI2BB2X1 U1349 ( .B0(n1571), .B1(n1917), .A0N(sigma6[1]), .A1N(n1931), .Y(
        n1746) );
  XOR2X1 U1350 ( .A(n1572), .B(L6_8[1]), .Y(n1571) );
  XOR2X1 U1351 ( .A(n1573), .B(n1574), .Y(n1572) );
  XOR2X1 U1352 ( .A(n1575), .B(n1576), .Y(n1574) );
  OAI2BB2X1 U1353 ( .B0(n1579), .B1(n1917), .A0N(sigma6[2]), .A1N(n1931), .Y(
        n1747) );
  XOR2X1 U1354 ( .A(n1580), .B(L6_8[2]), .Y(n1579) );
  XOR2X1 U1355 ( .A(n1581), .B(n1582), .Y(n1580) );
  XOR2X1 U1356 ( .A(n1583), .B(n1584), .Y(n1582) );
  OAI2BB2X1 U1357 ( .B0(n1651), .B1(n1905), .A0N(sigma6[11]), .A1N(n1927), .Y(
        n1756) );
  XOR2X1 U1358 ( .A(n1652), .B(L6_8[11]), .Y(n1651) );
  XOR2X1 U1359 ( .A(n1653), .B(n1654), .Y(n1652) );
  OAI2BB2X1 U1360 ( .B0(n1659), .B1(n1908), .A0N(sigma6[12]), .A1N(n1926), .Y(
        n1757) );
  XOR2X1 U1361 ( .A(n1660), .B(L6_8[12]), .Y(n1659) );
  XOR2X1 U1362 ( .A(n1661), .B(n1662), .Y(n1660) );
  XOR2X1 U1363 ( .A(n1663), .B(n1664), .Y(n1662) );
  OAI2BB2X1 U1364 ( .B0(n11), .B1(n1923), .A0N(sigma5[1]), .A1N(n1926), .Y(
        n1759) );
  XOR2X1 U1365 ( .A(n12), .B(L5_8[1]), .Y(n11) );
  XOR2X1 U1366 ( .A(n13), .B(n14), .Y(n12) );
  XOR2X1 U1367 ( .A(n15), .B(n16), .Y(n14) );
  OAI2BB2X1 U1368 ( .B0(n19), .B1(n1924), .A0N(sigma5[2]), .A1N(n1927), .Y(
        n1760) );
  XOR2X1 U1369 ( .A(n23), .B(n24), .Y(n22) );
  OAI2BB2X1 U1370 ( .B0(n155), .B1(n1921), .A0N(sigma4[6]), .A1N(n1930), .Y(
        n1777) );
  XOR2X1 U1371 ( .A(n156), .B(L4_8[6]), .Y(n155) );
  XOR2X1 U1372 ( .A(n157), .B(n158), .Y(n156) );
  OAI2BB2X1 U1373 ( .B0(n195), .B1(n1919), .A0N(sigma4[11]), .A1N(n1928), .Y(
        n1782) );
  XOR2X1 U1374 ( .A(n196), .B(L4_8[11]), .Y(n195) );
  XOR2X1 U1375 ( .A(n197), .B(n198), .Y(n196) );
  OAI2BB2X1 U1376 ( .B0(n299), .B1(n1920), .A0N(sigma3[11]), .A1N(n1944), .Y(
        n1795) );
  XOR2X1 U1377 ( .A(n300), .B(L3_8[11]), .Y(n299) );
  XOR2X1 U1378 ( .A(n301), .B(n302), .Y(n300) );
  OAI2BB2X1 U1379 ( .B0(n371), .B1(n1921), .A0N(sigma2[7]), .A1N(n1941), .Y(
        n1804) );
  XOR2X1 U1380 ( .A(n372), .B(L2_8[7]), .Y(n371) );
  XOR2X1 U1381 ( .A(n373), .B(n374), .Y(n372) );
  OAI2BB2X1 U1382 ( .B0(n531), .B1(n1924), .A0N(sigma16[1]), .A1N(n1935), .Y(
        n1824) );
  XOR2X1 U1383 ( .A(n532), .B(L16_8[1]), .Y(n531) );
  XOR2X1 U1384 ( .A(n533), .B(n534), .Y(n532) );
  XOR2X1 U1385 ( .A(n535), .B(n536), .Y(n534) );
  OAI2BB2X1 U1386 ( .B0(n563), .B1(n1905), .A0N(sigma16[5]), .A1N(n1940), .Y(
        n1828) );
  XOR2X1 U1387 ( .A(n564), .B(L16_8[5]), .Y(n563) );
  XOR2X1 U1388 ( .A(n565), .B(n566), .Y(n564) );
  XOR2X1 U1389 ( .A(n567), .B(n568), .Y(n566) );
  OAI2BB2X1 U1390 ( .B0(n587), .B1(n1905), .A0N(sigma16[8]), .A1N(n1935), .Y(
        n1831) );
  XOR2X1 U1391 ( .A(n588), .B(L16_8[8]), .Y(n587) );
  XOR2X1 U1392 ( .A(n589), .B(n590), .Y(n588) );
  XOR2X1 U1393 ( .A(n591), .B(n592), .Y(n590) );
  OAI2BB2X1 U1394 ( .B0(n643), .B1(n1906), .A0N(sigma14[2]), .A1N(n1936), .Y(
        n1838) );
  XOR2X1 U1395 ( .A(n644), .B(L14_8[2]), .Y(n643) );
  XOR2X1 U1396 ( .A(n645), .B(n646), .Y(n644) );
  OAI2BB2X1 U1397 ( .B0(n747), .B1(n1907), .A0N(sigma15[2]), .A1N(n1938), .Y(
        n1851) );
  XOR2X1 U1398 ( .A(n748), .B(L15_8[2]), .Y(n747) );
  XOR2X1 U1399 ( .A(n749), .B(n750), .Y(n748) );
  OAI2BB2X1 U1400 ( .B0(n851), .B1(n1908), .A0N(sigma13[2]), .A1N(n1940), .Y(
        n1864) );
  XOR2X1 U1401 ( .A(n852), .B(L13_8[2]), .Y(n851) );
  XOR2X1 U1402 ( .A(n853), .B(n854), .Y(n852) );
  OAI2BB2X1 U1403 ( .B0(n859), .B1(n1908), .A0N(sigma13[3]), .A1N(n1940), .Y(
        n1865) );
  XOR2X1 U1404 ( .A(n860), .B(L13_8[3]), .Y(n859) );
  XOR2X1 U1405 ( .A(n861), .B(n862), .Y(n860) );
  OAI2BB2X1 U1406 ( .B0(n883), .B1(n1909), .A0N(sigma13[6]), .A1N(n1940), .Y(
        n1868) );
  XOR2X1 U1407 ( .A(n884), .B(L13_8[6]), .Y(n883) );
  XOR2X1 U1408 ( .A(n885), .B(n886), .Y(n884) );
  OAI2BB2X1 U1409 ( .B0(n891), .B1(n1909), .A0N(sigma13[7]), .A1N(n1940), .Y(
        n1869) );
  XOR2X1 U1410 ( .A(n897), .B(n898), .Y(n893) );
  OAI2BB2X1 U1411 ( .B0(n923), .B1(n1909), .A0N(sigma13[11]), .A1N(n1941), .Y(
        n1873) );
  XOR2X1 U1412 ( .A(n924), .B(L13_8[11]), .Y(n923) );
  XOR2X1 U1413 ( .A(n925), .B(n926), .Y(n924) );
  OAI2BB2X1 U1414 ( .B0(n1547), .B1(n1917), .A0N(sigma7[11]), .A1N(n1933), .Y(
        n1743) );
  XOR2X1 U1415 ( .A(n1548), .B(L7_8[11]), .Y(n1547) );
  XOR2X1 U1416 ( .A(n1549), .B(n1550), .Y(n1548) );
  OAI2BB2X1 U1417 ( .B0(n1611), .B1(n1918), .A0N(sigma6[6]), .A1N(n1929), .Y(
        n1751) );
  XOR2X1 U1418 ( .A(n1612), .B(L6_8[6]), .Y(n1611) );
  XOR2X1 U1419 ( .A(n1613), .B(n1614), .Y(n1612) );
  OAI2BB2X1 U1420 ( .B0(n1539), .B1(n1917), .A0N(sigma7[10]), .A1N(n1933), .Y(
        n1742) );
  XOR2X1 U1421 ( .A(n1540), .B(L7_8[10]), .Y(n1539) );
  XOR2X1 U1422 ( .A(n1541), .B(n1542), .Y(n1540) );
  OAI2BB2X1 U1423 ( .B0(n1411), .B1(n1915), .A0N(sigma8[7]), .A1N(n1931), .Y(
        n1726) );
  XOR2X1 U1424 ( .A(n1412), .B(L8_8[7]), .Y(n1411) );
  XOR2X1 U1425 ( .A(n1413), .B(n1414), .Y(n1412) );
  XOR2X1 U1426 ( .A(n1417), .B(n1418), .Y(n1413) );
  OAI2BB2X1 U1427 ( .B0(n683), .B1(n1906), .A0N(sigma14[7]), .A1N(n1936), .Y(
        n1843) );
  XOR2X1 U1428 ( .A(n684), .B(L14_8[7]), .Y(n683) );
  XOR2X1 U1429 ( .A(n685), .B(n686), .Y(n684) );
  OAI2BB2X1 U1430 ( .B0(n811), .B1(n1908), .A0N(sigma15[10]), .A1N(n1939), .Y(
        n1859) );
  XOR2X1 U1431 ( .A(n812), .B(L15_8[10]), .Y(n811) );
  XOR2X1 U1432 ( .A(n813), .B(n814), .Y(n812) );
  OAI2BB2X1 U1433 ( .B0(n995), .B1(n1910), .A0N(sigma12[7]), .A1N(n1942), .Y(
        n1674) );
  XOR2X1 U1434 ( .A(n996), .B(L12_8[7]), .Y(n995) );
  XOR2X1 U1435 ( .A(n997), .B(n998), .Y(n996) );
  OAI2BB2X1 U1436 ( .B0(n779), .B1(n1907), .A0N(sigma15[6]), .A1N(n1938), .Y(
        n1855) );
  XOR2X1 U1437 ( .A(n780), .B(L15_8[6]), .Y(n779) );
  XOR2X1 U1438 ( .A(n781), .B(n782), .Y(n780) );
  OAI2BB2X1 U1439 ( .B0(n1523), .B1(n1917), .A0N(sigma7[8]), .A1N(n1934), .Y(
        n1740) );
  XOR2X1 U1440 ( .A(n1524), .B(L7_8[8]), .Y(n1523) );
  XOR2X1 U1441 ( .A(n1525), .B(n1526), .Y(n1524) );
  OAI2BB2X1 U1442 ( .B0(n1419), .B1(n1915), .A0N(sigma8[8]), .A1N(n1932), .Y(
        n1727) );
  XOR2X1 U1443 ( .A(n1420), .B(L8_8[8]), .Y(n1419) );
  XOR2X1 U1444 ( .A(n1422), .B(n1421), .Y(n1420) );
  OAI2BB2X1 U1445 ( .B0(n1507), .B1(n1917), .A0N(sigma7[6]), .A1N(n1934), .Y(
        n1738) );
  XOR2X1 U1446 ( .A(n1508), .B(L7_8[6]), .Y(n1507) );
  XOR2X1 U1447 ( .A(n1509), .B(n1510), .Y(n1508) );
  OAI2BB2X1 U1448 ( .B0(n1619), .B1(n1918), .A0N(sigma6[7]), .A1N(n1928), .Y(
        n1752) );
  XOR2X1 U1449 ( .A(n1620), .B(L6_8[7]), .Y(n1619) );
  XOR2X1 U1450 ( .A(n1621), .B(n1622), .Y(n1620) );
  OAI2BB2X1 U1451 ( .B0(n691), .B1(n1906), .A0N(sigma14[8]), .A1N(n1937), .Y(
        n1844) );
  XOR2X1 U1452 ( .A(n692), .B(L14_8[8]), .Y(n691) );
  XOR2X1 U1453 ( .A(n693), .B(n694), .Y(n692) );
  OAI2BB2X1 U1454 ( .B0(n1099), .B1(n1911), .A0N(sigma11[7]), .A1N(n1944), .Y(
        n1687) );
  XOR2X1 U1455 ( .A(n1100), .B(L11_8[7]), .Y(n1099) );
  XOR2X1 U1456 ( .A(n1101), .B(n1102), .Y(n1100) );
  XOR2X1 U1457 ( .A(n1105), .B(n1106), .Y(n1101) );
  OAI2BB2X1 U1458 ( .B0(n1643), .B1(n1918), .A0N(sigma6[10]), .A1N(n1927), .Y(
        n1755) );
  XOR2X1 U1459 ( .A(n1644), .B(L6_8[10]), .Y(n1643) );
  XOR2X1 U1460 ( .A(n1645), .B(n1646), .Y(n1644) );
  XOR2X1 U1461 ( .A(n1647), .B(n1648), .Y(n1646) );
  OAI2BB2X1 U1462 ( .B0(n1315), .B1(n1914), .A0N(sigma9[8]), .A1N(n1928), .Y(
        n1714) );
  XOR2X1 U1463 ( .A(n1316), .B(L9_8[8]), .Y(n1315) );
  XOR2X1 U1464 ( .A(n1317), .B(n1318), .Y(n1316) );
  OAI2BB2X1 U1465 ( .B0(n1123), .B1(n1912), .A0N(sigma11[10]), .A1N(n1945), 
        .Y(n1690) );
  XOR2X1 U1466 ( .A(n1124), .B(L11_8[10]), .Y(n1123) );
  XOR2X1 U1467 ( .A(n1125), .B(n1126), .Y(n1124) );
  OAI2BB2X1 U1468 ( .B0(n715), .B1(n1907), .A0N(sigma14[11]), .A1N(n1937), .Y(
        n1847) );
  XOR2X1 U1469 ( .A(n716), .B(L14_8[11]), .Y(n715) );
  XOR2X1 U1470 ( .A(n717), .B(n718), .Y(n716) );
  OAI2BB2X1 U1471 ( .B0(n899), .B1(n1909), .A0N(sigma13[8]), .A1N(n1941), .Y(
        n1870) );
  XOR2X1 U1472 ( .A(n900), .B(L13_8[8]), .Y(n899) );
  XOR2X1 U1473 ( .A(n901), .B(n902), .Y(n900) );
  XOR2X1 U1474 ( .A(n905), .B(n906), .Y(n901) );
  OAI2BB2X1 U1475 ( .B0(n987), .B1(n1910), .A0N(sigma12[6]), .A1N(n1942), .Y(
        n1673) );
  XOR2X1 U1476 ( .A(n988), .B(L12_8[6]), .Y(n987) );
  XOR2X1 U1477 ( .A(n989), .B(n990), .Y(n988) );
  OAI2BB2X1 U1478 ( .B0(n603), .B1(n1905), .A0N(sigma16[10]), .A1N(n1935), .Y(
        n1833) );
  XOR2X1 U1479 ( .A(n604), .B(L16_8[10]), .Y(n603) );
  XOR2X1 U1480 ( .A(n605), .B(n606), .Y(n604) );
  XOR2X1 U1481 ( .A(n609), .B(n610), .Y(n605) );
  OAI2BB2X1 U1482 ( .B0(n1403), .B1(n1915), .A0N(sigma8[6]), .A1N(n1931), .Y(
        n1725) );
  XOR2X1 U1483 ( .A(n1404), .B(L8_8[6]), .Y(n1403) );
  XOR2X1 U1484 ( .A(n1405), .B(n1406), .Y(n1404) );
  OAI2BB2X1 U1485 ( .B0(n1339), .B1(n1914), .A0N(sigma9[11]), .A1N(n1929), .Y(
        n1717) );
  XOR2X1 U1486 ( .A(n1340), .B(L9_8[11]), .Y(n1339) );
  XOR2X1 U1487 ( .A(n1341), .B(n1342), .Y(n1340) );
  OAI2BB2X1 U1488 ( .B0(n1083), .B1(n1911), .A0N(sigma11[5]), .A1N(n1944), .Y(
        n1685) );
  XOR2X1 U1489 ( .A(n1084), .B(L11_8[5]), .Y(n1083) );
  XOR2X1 U1490 ( .A(n1085), .B(n1086), .Y(n1084) );
  XOR2X1 U1491 ( .A(n1089), .B(n1090), .Y(n1085) );
  OAI2BB2X1 U1492 ( .B0(n1003), .B1(n1910), .A0N(sigma12[8]), .A1N(n1943), .Y(
        n1675) );
  XOR2X1 U1493 ( .A(n1004), .B(L12_8[8]), .Y(n1003) );
  XOR2X1 U1494 ( .A(n1005), .B(n1006), .Y(n1004) );
  OAI2BB2X1 U1495 ( .B0(n1299), .B1(n1914), .A0N(sigma9[6]), .A1N(n1929), .Y(
        n1712) );
  XOR2X1 U1496 ( .A(n1300), .B(L9_8[6]), .Y(n1299) );
  XOR2X1 U1497 ( .A(n1301), .B(n1302), .Y(n1300) );
  OAI2BB2X1 U1498 ( .B0(n1235), .B1(n1913), .A0N(sigma10[11]), .A1N(n1926), 
        .Y(n1704) );
  XOR2X1 U1499 ( .A(n1236), .B(L10_8[11]), .Y(n1235) );
  XOR2X1 U1500 ( .A(n1237), .B(n1238), .Y(n1236) );
  OAI2BB2X1 U1501 ( .B0(n1011), .B1(n1910), .A0N(sigma12[9]), .A1N(n1943), .Y(
        n1676) );
  XOR2X1 U1502 ( .A(n1012), .B(L12_8[9]), .Y(n1011) );
  XOR2X1 U1503 ( .A(n1013), .B(n1014), .Y(n1012) );
  OAI2BB2X1 U1504 ( .B0(n1195), .B1(n1913), .A0N(sigma10[6]), .A1N(n1925), .Y(
        n1699) );
  XOR2X1 U1505 ( .A(n1196), .B(L10_8[6]), .Y(n1195) );
  XOR2X1 U1506 ( .A(n1197), .B(n1198), .Y(n1196) );
  OAI2BB2X1 U1507 ( .B0(n579), .B1(n1905), .A0N(sigma16[7]), .A1N(n1935), .Y(
        n1830) );
  XOR2X1 U1508 ( .A(n580), .B(L16_8[7]), .Y(n579) );
  XOR2X1 U1509 ( .A(n581), .B(n582), .Y(n580) );
  XOR2X1 U1510 ( .A(n583), .B(n584), .Y(n582) );
  OAI2BB2X1 U1511 ( .B0(n1115), .B1(n1912), .A0N(sigma11[9]), .A1N(n1945), .Y(
        n1689) );
  XOR2X1 U1512 ( .A(n1121), .B(n1122), .Y(n1117) );
  OAI2BB2X1 U1513 ( .B0(n59), .B1(n1924), .A0N(sigma5[7]), .A1N(n1932), .Y(
        n1765) );
  XOR2X1 U1514 ( .A(n60), .B(L5_8[7]), .Y(n59) );
  XOR2X1 U1515 ( .A(n61), .B(n62), .Y(n60) );
  OAI2BB2X1 U1516 ( .B0(n51), .B1(n1925), .A0N(sigma5[6]), .A1N(n1931), .Y(
        n1764) );
  XOR2X1 U1517 ( .A(n52), .B(L5_8[6]), .Y(n51) );
  XOR2X1 U1518 ( .A(n53), .B(n54), .Y(n52) );
  OAI2BB2X1 U1519 ( .B0(n819), .B1(n1908), .A0N(sigma15[11]), .A1N(n1939), .Y(
        n1860) );
  XOR2X1 U1520 ( .A(n820), .B(L15_8[11]), .Y(n819) );
  XOR2X1 U1521 ( .A(n821), .B(n822), .Y(n820) );
  OAI2BB2X1 U1522 ( .B0(n907), .B1(n1909), .A0N(sigma13[9]), .A1N(n1941), .Y(
        n1871) );
  XOR2X1 U1523 ( .A(n908), .B(L13_8[9]), .Y(n907) );
  XOR2X1 U1524 ( .A(n909), .B(n910), .Y(n908) );
  OAI2BB2X1 U1525 ( .B0(n699), .B1(n1906), .A0N(sigma14[9]), .A1N(n1937), .Y(
        n1845) );
  XOR2X1 U1526 ( .A(n700), .B(L14_8[9]), .Y(n699) );
  XOR2X1 U1527 ( .A(n701), .B(n702), .Y(n700) );
  OAI2BB2X1 U1528 ( .B0(n1443), .B1(n1916), .A0N(sigma8[11]), .A1N(n1932), .Y(
        n1730) );
  XOR2X1 U1529 ( .A(n1444), .B(L8_8[11]), .Y(n1443) );
  XOR2X1 U1530 ( .A(n1445), .B(n1446), .Y(n1444) );
  OAI2BB2X1 U1531 ( .B0(n1587), .B1(n1918), .A0N(sigma6[3]), .A1N(n1930), .Y(
        n1748) );
  XOR2X1 U1532 ( .A(n1588), .B(L6_8[3]), .Y(n1587) );
  XOR2X1 U1533 ( .A(n1589), .B(n1590), .Y(n1588) );
  OAI2BB2X1 U1534 ( .B0(n1531), .B1(n1917), .A0N(sigma7[9]), .A1N(n1934), .Y(
        n1741) );
  XOR2X1 U1535 ( .A(n1532), .B(L7_8[9]), .Y(n1531) );
  XOR2X1 U1536 ( .A(n1533), .B(n1534), .Y(n1532) );
  OAI2BB2X1 U1537 ( .B0(n1515), .B1(n1917), .A0N(sigma7[7]), .A1N(n1934), .Y(
        n1739) );
  XOR2X1 U1538 ( .A(n1516), .B(L7_8[7]), .Y(n1515) );
  XOR2X1 U1539 ( .A(n1517), .B(n1518), .Y(n1516) );
  OAI2BB2X1 U1540 ( .B0(n1379), .B1(n1915), .A0N(sigma8[3]), .A1N(n1930), .Y(
        n1722) );
  XOR2X1 U1541 ( .A(n1380), .B(L8_8[3]), .Y(n1379) );
  XOR2X1 U1542 ( .A(n1381), .B(n1382), .Y(n1380) );
  OAI2BB2X1 U1543 ( .B0(n163), .B1(n1920), .A0N(sigma4[7]), .A1N(n1930), .Y(
        n1778) );
  XOR2X1 U1544 ( .A(n164), .B(L4_8[7]), .Y(n163) );
  XOR2X1 U1545 ( .A(n165), .B(n166), .Y(n164) );
  OAI2BB2X1 U1546 ( .B0(n1267), .B1(n1914), .A0N(sigma9[2]), .A1N(n1928), .Y(
        n1708) );
  XOR2X1 U1547 ( .A(n1268), .B(L9_8[2]), .Y(n1267) );
  XOR2X1 U1548 ( .A(n1269), .B(n1270), .Y(n1268) );
  OAI2BB2X1 U1549 ( .B0(n755), .B1(n1907), .A0N(sigma15[3]), .A1N(n1938), .Y(
        n1852) );
  XOR2X1 U1550 ( .A(n756), .B(L15_8[3]), .Y(n755) );
  XOR2X1 U1551 ( .A(n757), .B(n758), .Y(n756) );
  OAI2BB2X1 U1552 ( .B0(n67), .B1(n1923), .A0N(sigma5[8]), .A1N(n1933), .Y(
        n1766) );
  XOR2X1 U1553 ( .A(n68), .B(L5_8[8]), .Y(n67) );
  XOR2X1 U1554 ( .A(n69), .B(n70), .Y(n68) );
  OAI2BB2X1 U1555 ( .B0(n75), .B1(n1923), .A0N(sigma5[9]), .A1N(n1926), .Y(
        n1767) );
  XOR2X1 U1556 ( .A(n76), .B(L5_8[9]), .Y(n75) );
  XOR2X1 U1557 ( .A(n77), .B(n78), .Y(n76) );
  OAI2BB2X1 U1558 ( .B0(n187), .B1(n1920), .A0N(sigma4[10]), .A1N(n1928), .Y(
        n1781) );
  XOR2X1 U1559 ( .A(n188), .B(L4_8[10]), .Y(n187) );
  XOR2X1 U1560 ( .A(n189), .B(n190), .Y(n188) );
  XOR2X1 U1561 ( .A(n191), .B(n192), .Y(n190) );
  OAI2BB2X1 U1562 ( .B0(n1219), .B1(n1913), .A0N(sigma10[9]), .A1N(n1925), .Y(
        n1702) );
  XOR2X1 U1563 ( .A(n1220), .B(L10_8[9]), .Y(n1219) );
  XOR2X1 U1564 ( .A(n1221), .B(n1222), .Y(n1220) );
  OAI2BB2X1 U1565 ( .B0(n83), .B1(n1923), .A0N(sigma5[10]), .A1N(n1934), .Y(
        n1768) );
  XOR2X1 U1566 ( .A(n84), .B(L5_8[10]), .Y(n83) );
  XOR2X1 U1567 ( .A(n85), .B(n86), .Y(n84) );
  OAI2BB2X1 U1568 ( .B0(n123), .B1(n1922), .A0N(sigma4[2]), .A1N(n1932), .Y(
        n1773) );
  XOR2X1 U1569 ( .A(n124), .B(L4_8[2]), .Y(n123) );
  XOR2X1 U1570 ( .A(n125), .B(n126), .Y(n124) );
  OAI2BB2X1 U1571 ( .B0(n955), .B1(n1910), .A0N(sigma12[2]), .A1N(n1942), .Y(
        n1669) );
  XOR2X1 U1572 ( .A(n956), .B(L12_8[2]), .Y(n955) );
  XOR2X1 U1573 ( .A(n957), .B(n958), .Y(n956) );
  XOR2X1 U1574 ( .A(n959), .B(n960), .Y(n958) );
  OAI2BB2X1 U1575 ( .B0(n1131), .B1(n1912), .A0N(sigma11[11]), .A1N(n1945), 
        .Y(n1691) );
  XOR2X1 U1576 ( .A(n1132), .B(L11_8[11]), .Y(n1131) );
  XOR2X1 U1577 ( .A(n1133), .B(n1134), .Y(n1132) );
  XOR2X1 U1578 ( .A(n1137), .B(n1138), .Y(n1133) );
  OAI2BB2X1 U1579 ( .B0(n1163), .B1(n1912), .A0N(sigma10[2]), .A1N(n1946), .Y(
        n1695) );
  XOR2X1 U1580 ( .A(n1164), .B(L10_8[2]), .Y(n1163) );
  XOR2X1 U1581 ( .A(n1165), .B(n1166), .Y(n1164) );
  XOR2X1 U1582 ( .A(n1167), .B(n1168), .Y(n1166) );
  OAI2BB2X1 U1583 ( .B0(n1227), .B1(n1913), .A0N(sigma10[10]), .A1N(n1927), 
        .Y(n1703) );
  XOR2X1 U1584 ( .A(n1228), .B(L10_8[10]), .Y(n1227) );
  XOR2X1 U1585 ( .A(n1229), .B(n1230), .Y(n1228) );
  OAI2BB2X1 U1586 ( .B0(n1275), .B1(n1914), .A0N(sigma9[3]), .A1N(n1928), .Y(
        n1709) );
  XOR2X1 U1587 ( .A(n1276), .B(L9_8[3]), .Y(n1275) );
  XOR2X1 U1588 ( .A(n1277), .B(n1278), .Y(n1276) );
  OAI2BB2X1 U1589 ( .B0(n1467), .B1(n1916), .A0N(sigma7[1]), .A1N(n1933), .Y(
        n1733) );
  XOR2X1 U1590 ( .A(n1468), .B(L7_8[1]), .Y(n1467) );
  XOR2X1 U1591 ( .A(n1469), .B(n1470), .Y(n1468) );
  OAI2BB2X1 U1592 ( .B0(n1483), .B1(n1916), .A0N(sigma7[3]), .A1N(n1933), .Y(
        n1735) );
  XOR2X1 U1593 ( .A(n1484), .B(L7_8[3]), .Y(n1483) );
  XOR2X1 U1594 ( .A(n1485), .B(n1486), .Y(n1484) );
  OAI2BB2X1 U1595 ( .B0(n27), .B1(n1925), .A0N(sigma5[3]), .A1N(n1929), .Y(
        n1761) );
  XOR2X1 U1596 ( .A(n28), .B(L5_8[3]), .Y(n27) );
  XOR2X1 U1597 ( .A(n29), .B(n30), .Y(n28) );
  OAI2BB2X1 U1598 ( .B0(n227), .B1(n1919), .A0N(sigma3[2]), .A1N(n1926), .Y(
        n1786) );
  XOR2X1 U1599 ( .A(n228), .B(L3_8[2]), .Y(n227) );
  XOR2X1 U1600 ( .A(n229), .B(n230), .Y(n228) );
  OAI2BB2X1 U1601 ( .B0(n235), .B1(n1919), .A0N(sigma3[3]), .A1N(n1926), .Y(
        n1787) );
  XOR2X1 U1602 ( .A(n236), .B(L3_8[3]), .Y(n235) );
  XOR2X1 U1603 ( .A(n237), .B(n238), .Y(n236) );
  OAI2BB2X1 U1604 ( .B0(n267), .B1(n1919), .A0N(sigma3[7]), .A1N(n1945), .Y(
        n1791) );
  XOR2X1 U1605 ( .A(n271), .B(n272), .Y(n270) );
  OAI2BB2X1 U1606 ( .B0(n275), .B1(n1923), .A0N(sigma3[8]), .A1N(n1945), .Y(
        n1792) );
  XOR2X1 U1607 ( .A(n276), .B(L3_8[8]), .Y(n275) );
  XOR2X1 U1608 ( .A(n277), .B(n278), .Y(n276) );
  OAI2BB2X1 U1609 ( .B0(n283), .B1(n1919), .A0N(sigma3[9]), .A1N(n1944), .Y(
        n1793) );
  XOR2X1 U1610 ( .A(n284), .B(L3_8[9]), .Y(n283) );
  XOR2X1 U1611 ( .A(n285), .B(n286), .Y(n284) );
  OAI2BB2X1 U1612 ( .B0(n291), .B1(n1920), .A0N(sigma3[10]), .A1N(n1944), .Y(
        n1794) );
  XOR2X1 U1613 ( .A(n292), .B(L3_8[10]), .Y(n291) );
  XOR2X1 U1614 ( .A(n293), .B(n294), .Y(n292) );
  OAI2BB2X1 U1615 ( .B0(n315), .B1(n1920), .A0N(sigma2[0]), .A1N(n1943), .Y(
        n1797) );
  XOR2X1 U1616 ( .A(n316), .B(L2_8[0]), .Y(n315) );
  XOR2X1 U1617 ( .A(n317), .B(n318), .Y(n316) );
  XOR2X1 U1618 ( .A(n319), .B(n320), .Y(n318) );
  OAI2BB2X1 U1619 ( .B0(n323), .B1(n1920), .A0N(sigma2[1]), .A1N(n1943), .Y(
        n1798) );
  XOR2X1 U1620 ( .A(n324), .B(L2_8[1]), .Y(n323) );
  XOR2X1 U1621 ( .A(n325), .B(n326), .Y(n324) );
  OAI2BB2X1 U1622 ( .B0(n331), .B1(n1920), .A0N(sigma2[2]), .A1N(n1943), .Y(
        n1799) );
  XOR2X1 U1623 ( .A(n332), .B(L2_8[2]), .Y(n331) );
  XOR2X1 U1624 ( .A(n333), .B(n334), .Y(n332) );
  XOR2X1 U1625 ( .A(n335), .B(n336), .Y(n334) );
  OAI2BB2X1 U1626 ( .B0(n339), .B1(n1921), .A0N(sigma2[3]), .A1N(n1942), .Y(
        n1800) );
  XOR2X1 U1627 ( .A(n340), .B(L2_8[3]), .Y(n339) );
  XOR2X1 U1628 ( .A(n341), .B(n342), .Y(n340) );
  OAI2BB2X1 U1629 ( .B0(n379), .B1(n1921), .A0N(sigma2[8]), .A1N(n1941), .Y(
        n1805) );
  XOR2X1 U1630 ( .A(n380), .B(L2_8[8]), .Y(n379) );
  XOR2X1 U1631 ( .A(n381), .B(n382), .Y(n380) );
  OAI2BB2X1 U1632 ( .B0(n387), .B1(n1922), .A0N(sigma2[9]), .A1N(n1941), .Y(
        n1806) );
  XOR2X1 U1633 ( .A(n388), .B(L2_8[9]), .Y(n387) );
  XOR2X1 U1634 ( .A(n389), .B(n390), .Y(n388) );
  OAI2BB2X1 U1635 ( .B0(n395), .B1(n1922), .A0N(sigma2[10]), .A1N(n1940), .Y(
        n1807) );
  XOR2X1 U1636 ( .A(n399), .B(n400), .Y(n398) );
  OAI2BB2X1 U1637 ( .B0(n403), .B1(n1922), .A0N(sigma2[11]), .A1N(n1940), .Y(
        n1808) );
  XOR2X1 U1638 ( .A(n407), .B(n408), .Y(n406) );
  OAI2BB2X1 U1639 ( .B0(n435), .B1(n1923), .A0N(sigma1[2]), .A1N(n1939), .Y(
        n1812) );
  XOR2X1 U1640 ( .A(n439), .B(n440), .Y(n438) );
  OAI2BB2X1 U1641 ( .B0(n443), .B1(n1923), .A0N(sigma1[3]), .A1N(n1938), .Y(
        n1813) );
  XOR2X1 U1642 ( .A(n449), .B(n450), .Y(n445) );
  OAI2BB2X1 U1643 ( .B0(n467), .B1(n1924), .A0N(sigma1[6]), .A1N(n1937), .Y(
        n1816) );
  XOR2X1 U1644 ( .A(n468), .B(L1_8[6]), .Y(n467) );
  XOR2X1 U1645 ( .A(n469), .B(n470), .Y(n468) );
  OAI2BB2X1 U1646 ( .B0(n475), .B1(n1924), .A0N(sigma1[7]), .A1N(n1937), .Y(
        n1817) );
  XOR2X1 U1647 ( .A(n479), .B(n480), .Y(n478) );
  OAI2BB2X1 U1648 ( .B0(n483), .B1(n1924), .A0N(sigma1[8]), .A1N(n1937), .Y(
        n1818) );
  XOR2X1 U1649 ( .A(n484), .B(L1_8[8]), .Y(n483) );
  XOR2X1 U1650 ( .A(n485), .B(n486), .Y(n484) );
  OAI2BB2X1 U1651 ( .B0(n491), .B1(n1924), .A0N(sigma1[9]), .A1N(n1937), .Y(
        n1819) );
  XOR2X1 U1652 ( .A(n492), .B(L1_8[9]), .Y(n491) );
  XOR2X1 U1653 ( .A(n493), .B(n494), .Y(n492) );
  OAI2BB2X1 U1654 ( .B0(n499), .B1(n1925), .A0N(sigma1[10]), .A1N(n1936), .Y(
        n1820) );
  XOR2X1 U1655 ( .A(n500), .B(L1_8[10]), .Y(n499) );
  XOR2X1 U1656 ( .A(n501), .B(n502), .Y(n500) );
  OAI2BB2X1 U1657 ( .B0(n507), .B1(n1925), .A0N(sigma1[11]), .A1N(n1936), .Y(
        n1821) );
  XOR2X1 U1658 ( .A(n508), .B(L1_8[11]), .Y(n507) );
  XOR2X1 U1659 ( .A(n509), .B(n510), .Y(n508) );
  XOR2X1 U1660 ( .A(n511), .B(n512), .Y(n510) );
  OAI2BB2X1 U1661 ( .B0(n515), .B1(n1925), .A0N(sigma1[12]), .A1N(n1936), .Y(
        n1822) );
  XOR2X1 U1662 ( .A(n519), .B(n520), .Y(n518) );
  OAI2BB2X1 U1663 ( .B0(n547), .B1(n1924), .A0N(sigma16[3]), .A1N(n1934), .Y(
        n1826) );
  XOR2X1 U1664 ( .A(n548), .B(L16_8[3]), .Y(n547) );
  XOR2X1 U1665 ( .A(n549), .B(n550), .Y(n548) );
  XOR2X1 U1666 ( .A(n553), .B(n554), .Y(n549) );
  OAI2BB2X1 U1667 ( .B0(n635), .B1(n1906), .A0N(sigma14[1]), .A1N(n1936), .Y(
        n1837) );
  XOR2X1 U1668 ( .A(n636), .B(L14_8[1]), .Y(n635) );
  XOR2X1 U1669 ( .A(n637), .B(n638), .Y(n636) );
  OAI2BB2X1 U1670 ( .B0(n843), .B1(n1908), .A0N(sigma13[1]), .A1N(n1939), .Y(
        n1863) );
  XOR2X1 U1671 ( .A(n844), .B(L13_8[1]), .Y(n843) );
  XOR2X1 U1672 ( .A(n845), .B(n846), .Y(n844) );
  XNOR2X1 U1673 ( .A(L10_2[3]), .B(L10_1[3]), .Y(n1176) );
  XOR2X1 U1674 ( .A(L6_4[3]), .B(L6_3[3]), .Y(n1902) );
  XNOR2X1 U1675 ( .A(L15_2[3]), .B(L15_1[3]), .Y(n760) );
  OAI2BB2X1 U1676 ( .B0(n1251), .B1(n1913), .A0N(sigma9[0]), .A1N(n1928), .Y(
        n1706) );
  XOR2X1 U1677 ( .A(n1252), .B(L9_8[0]), .Y(n1251) );
  XOR2X1 U1678 ( .A(n1253), .B(n1254), .Y(n1252) );
  XOR2X1 U1679 ( .A(n1255), .B(n1256), .Y(n1254) );
  OAI2BB2X1 U1680 ( .B0(n1291), .B1(n1914), .A0N(sigma9[5]), .A1N(n1927), .Y(
        n1711) );
  XOR2X1 U1681 ( .A(n1292), .B(L9_8[5]), .Y(n1291) );
  XOR2X1 U1682 ( .A(n1293), .B(n1294), .Y(n1292) );
  XOR2X1 U1683 ( .A(n1297), .B(n1298), .Y(n1293) );
  OAI2BB2X1 U1684 ( .B0(n979), .B1(n1910), .A0N(sigma12[5]), .A1N(n1942), .Y(
        n1672) );
  XOR2X1 U1685 ( .A(n980), .B(L12_8[5]), .Y(n979) );
  XOR2X1 U1686 ( .A(n981), .B(n982), .Y(n980) );
  XOR2X1 U1687 ( .A(n985), .B(n986), .Y(n981) );
  OAI2BB2X1 U1688 ( .B0(n619), .B1(n1905), .A0N(sigma16[12]), .A1N(n1935), .Y(
        n1835) );
  XOR2X1 U1689 ( .A(n620), .B(L16_8[12]), .Y(n619) );
  XOR2X1 U1690 ( .A(n621), .B(n622), .Y(n620) );
  XOR2X1 U1691 ( .A(n623), .B(n624), .Y(n622) );
  OAI2BB2X1 U1692 ( .B0(n259), .B1(n1919), .A0N(sigma3[6]), .A1N(n1945), .Y(
        n1790) );
  XOR2X1 U1693 ( .A(n260), .B(L3_8[6]), .Y(n259) );
  XOR2X1 U1694 ( .A(n261), .B(n262), .Y(n260) );
  XOR2X1 U1695 ( .A(n263), .B(n264), .Y(n262) );
  XOR2X1 U1696 ( .A(n737), .B(n738), .Y(n733) );
  XOR2X1 U1697 ( .A(n873), .B(n874), .Y(n869) );
  OAI2BB2X1 U1698 ( .B0(n1139), .B1(n1912), .A0N(sigma11[12]), .A1N(n1945), 
        .Y(n1692) );
  XOR2X1 U1699 ( .A(n1140), .B(L11_8[12]), .Y(n1139) );
  XOR2X1 U1700 ( .A(n1141), .B(n1142), .Y(n1140) );
  XOR2X1 U1701 ( .A(n1145), .B(n1146), .Y(n1141) );
  OAI2BB2X1 U1702 ( .B0(n1563), .B1(n1917), .A0N(sigma6[0]), .A1N(n1932), .Y(
        n1745) );
  XOR2X1 U1703 ( .A(n1564), .B(L6_8[0]), .Y(n1563) );
  XOR2X1 U1704 ( .A(n1565), .B(n1566), .Y(n1564) );
  XOR2X1 U1705 ( .A(n1567), .B(n1568), .Y(n1566) );
  OAI2BB2X1 U1706 ( .B0(n107), .B1(n1922), .A0N(sigma4[0]), .A1N(n1933), .Y(
        n1771) );
  XOR2X1 U1707 ( .A(n108), .B(L4_8[0]), .Y(n107) );
  XOR2X1 U1708 ( .A(n109), .B(n110), .Y(n108) );
  XOR2X1 U1709 ( .A(n111), .B(n112), .Y(n110) );
  OAI2BB2X1 U1710 ( .B0(n203), .B1(n1919), .A0N(sigma4[12]), .A1N(n1927), .Y(
        n1783) );
  XOR2X1 U1711 ( .A(n204), .B(L4_8[12]), .Y(n203) );
  XOR2X1 U1712 ( .A(n205), .B(n206), .Y(n204) );
  XOR2X1 U1713 ( .A(n207), .B(n208), .Y(n206) );
  OAI2BB2X1 U1714 ( .B0(n827), .B1(n1918), .A0N(sigma15[12]), .A1N(n1939), .Y(
        n1861) );
  XOR2X1 U1715 ( .A(n828), .B(L15_8[12]), .Y(n827) );
  XOR2X1 U1716 ( .A(n829), .B(n830), .Y(n828) );
  XOR2X1 U1717 ( .A(n833), .B(n834), .Y(n829) );
  OAI2BB2X1 U1718 ( .B0(n211), .B1(n1919), .A0N(sigma3[0]), .A1N(n1926), .Y(
        n1784) );
  XOR2X1 U1719 ( .A(n212), .B(L3_8[0]), .Y(n211) );
  XOR2X1 U1720 ( .A(n213), .B(n214), .Y(n212) );
  XOR2X1 U1721 ( .A(n215), .B(n216), .Y(n214) );
  OAI2BB2X1 U1722 ( .B0(n1459), .B1(n1916), .A0N(sigma7[0]), .A1N(n1933), .Y(
        n1732) );
  XOR2X1 U1723 ( .A(n1460), .B(L7_8[0]), .Y(n1459) );
  XOR2X1 U1724 ( .A(n1461), .B(n1462), .Y(n1460) );
  XOR2X1 U1725 ( .A(n1463), .B(n1464), .Y(n1462) );
  OAI2BB2X1 U1726 ( .B0(n875), .B1(n1909), .A0N(sigma13[5]), .A1N(n1940), .Y(
        n1867) );
  XOR2X1 U1727 ( .A(n876), .B(L13_8[5]), .Y(n875) );
  XOR2X1 U1728 ( .A(n877), .B(n878), .Y(n876) );
  XOR2X1 U1729 ( .A(n881), .B(n882), .Y(n877) );
  OAI2BB2X1 U1730 ( .B0(n1347), .B1(n1915), .A0N(sigma9[12]), .A1N(n1930), .Y(
        n1718) );
  XOR2X1 U1731 ( .A(n1348), .B(L9_8[12]), .Y(n1347) );
  XOR2X1 U1732 ( .A(n1349), .B(n1350), .Y(n1348) );
  XOR2X1 U1733 ( .A(n1351), .B(n1352), .Y(n1350) );
  OAI2BB2X1 U1734 ( .B0(n147), .B1(n1921), .A0N(sigma4[5]), .A1N(n1930), .Y(
        n1776) );
  XOR2X1 U1735 ( .A(n148), .B(L4_8[5]), .Y(n147) );
  XOR2X1 U1736 ( .A(n149), .B(n150), .Y(n148) );
  XOR2X1 U1737 ( .A(n151), .B(n152), .Y(n150) );
  OAI2BB2X1 U1738 ( .B0(n931), .B1(n1909), .A0N(sigma13[12]), .A1N(n1941), .Y(
        n1874) );
  XOR2X1 U1739 ( .A(n932), .B(L13_8[12]), .Y(n931) );
  XOR2X1 U1740 ( .A(n933), .B(n934), .Y(n932) );
  XOR2X1 U1741 ( .A(n937), .B(n938), .Y(n933) );
  OAI2BB2X1 U1742 ( .B0(n1555), .B1(n1917), .A0N(sigma7[12]), .A1N(n1932), .Y(
        n1744) );
  XOR2X1 U1743 ( .A(n1556), .B(L7_8[12]), .Y(n1555) );
  XOR2X1 U1744 ( .A(n1557), .B(n1558), .Y(n1556) );
  XOR2X1 U1745 ( .A(n1559), .B(n1560), .Y(n1558) );
  OAI2BB2X1 U1746 ( .B0(n1355), .B1(n1915), .A0N(sigma8[0]), .A1N(n1930), .Y(
        n1719) );
  XOR2X1 U1747 ( .A(n1356), .B(L8_8[0]), .Y(n1355) );
  XOR2X1 U1748 ( .A(n1357), .B(n1358), .Y(n1356) );
  XOR2X1 U1749 ( .A(n1359), .B(n1360), .Y(n1358) );
  OAI2BB2X1 U1750 ( .B0(n1451), .B1(n1916), .A0N(sigma8[12]), .A1N(n1932), .Y(
        n1731) );
  XOR2X1 U1751 ( .A(n1452), .B(L8_8[12]), .Y(n1451) );
  XOR2X1 U1752 ( .A(n1453), .B(n1454), .Y(n1452) );
  XOR2X1 U1753 ( .A(n1457), .B(n1458), .Y(n1453) );
  OAI2BB2X1 U1754 ( .B0(n307), .B1(n1920), .A0N(sigma3[12]), .A1N(n1944), .Y(
        n1796) );
  XOR2X1 U1755 ( .A(n308), .B(L3_8[12]), .Y(n307) );
  XOR2X1 U1756 ( .A(n309), .B(n310), .Y(n308) );
  XOR2X1 U1757 ( .A(n311), .B(n312), .Y(n310) );
  OAI2BB2X1 U1758 ( .B0(n411), .B1(n1922), .A0N(sigma2[12]), .A1N(n1940), .Y(
        n1809) );
  XOR2X1 U1759 ( .A(n412), .B(L2_8[12]), .Y(n411) );
  XOR2X1 U1760 ( .A(n413), .B(n414), .Y(n412) );
  XOR2X1 U1761 ( .A(n415), .B(n416), .Y(n414) );
  OAI2BB2X1 U1762 ( .B0(n1019), .B1(n1910), .A0N(sigma12[10]), .A1N(n1943), 
        .Y(n1677) );
  XOR2X1 U1763 ( .A(n1020), .B(L12_8[10]), .Y(n1019) );
  XOR2X1 U1764 ( .A(n1021), .B(n1022), .Y(n1020) );
  XOR2X1 U1765 ( .A(n1025), .B(n1026), .Y(n1021) );
  OAI2BB2X1 U1766 ( .B0(n171), .B1(n1920), .A0N(sigma4[8]), .A1N(n1929), .Y(
        n1779) );
  XOR2X1 U1767 ( .A(n172), .B(L4_8[8]), .Y(n171) );
  XOR2X1 U1768 ( .A(n173), .B(n174), .Y(n172) );
  OAI2BB2X1 U1769 ( .B0(n739), .B1(n1907), .A0N(sigma15[1]), .A1N(n1938), .Y(
        n1850) );
  XOR2X1 U1770 ( .A(n740), .B(L15_8[1]), .Y(n739) );
  XOR2X1 U1771 ( .A(n741), .B(n742), .Y(n740) );
  OAI2BB2X1 U1772 ( .B0(n803), .B1(n1908), .A0N(sigma15[9]), .A1N(n1939), .Y(
        n1858) );
  XOR2X1 U1773 ( .A(n804), .B(L15_8[9]), .Y(n803) );
  XOR2X1 U1774 ( .A(n805), .B(n806), .Y(n804) );
  OAI2BB2X1 U1775 ( .B0(n131), .B1(n1921), .A0N(sigma4[3]), .A1N(n1931), .Y(
        n1774) );
  XOR2X1 U1776 ( .A(n132), .B(L4_8[3]), .Y(n131) );
  XOR2X1 U1777 ( .A(n133), .B(n134), .Y(n132) );
  OAI2BB2X1 U1778 ( .B0(n179), .B1(n1920), .A0N(sigma4[9]), .A1N(n1928), .Y(
        n1780) );
  XOR2X1 U1779 ( .A(n180), .B(L4_8[9]), .Y(n179) );
  XOR2X1 U1780 ( .A(n181), .B(n182), .Y(n180) );
  OAI2BB2X1 U1781 ( .B0(n1427), .B1(n1916), .A0N(sigma8[9]), .A1N(n1932), .Y(
        n1728) );
  XOR2X1 U1782 ( .A(n1428), .B(L8_8[9]), .Y(n1427) );
  XOR2X1 U1783 ( .A(n1429), .B(n1430), .Y(n1428) );
  OAI2BB2X1 U1784 ( .B0(n219), .B1(n1919), .A0N(sigma3[1]), .A1N(n1927), .Y(
        n1785) );
  XOR2X1 U1785 ( .A(n220), .B(L3_8[1]), .Y(n219) );
  XOR2X1 U1786 ( .A(n221), .B(n222), .Y(n220) );
  OAI2BB2X1 U1787 ( .B0(n1395), .B1(n1915), .A0N(sigma8[5]), .A1N(n1931), .Y(
        n1724) );
  XOR2X1 U1788 ( .A(n1396), .B(L8_8[5]), .Y(n1395) );
  XOR2X1 U1789 ( .A(n1397), .B(n1398), .Y(n1396) );
  OAI2BB2X1 U1790 ( .B0(n763), .B1(n1907), .A0N(sigma15[4]), .A1N(n1938), .Y(
        n1853) );
  XOR2X1 U1791 ( .A(n764), .B(L15_8[4]), .Y(n763) );
  XOR2X1 U1792 ( .A(n765), .B(n766), .Y(n764) );
  OAI2BB2X1 U1793 ( .B0(n1147), .B1(n1912), .A0N(sigma10[0]), .A1N(n1945), .Y(
        n1693) );
  XOR2X1 U1794 ( .A(n1148), .B(L10_8[0]), .Y(n1147) );
  XOR2X1 U1795 ( .A(n1149), .B(n1150), .Y(n1148) );
  OAI2BB2X1 U1796 ( .B0(n835), .B1(n1908), .A0N(sigma13[0]), .A1N(n1939), .Y(
        n1862) );
  XOR2X1 U1797 ( .A(n836), .B(L13_8[0]), .Y(n835) );
  XOR2X1 U1798 ( .A(n837), .B(n838), .Y(n836) );
  OAI2BB2X1 U1799 ( .B0(n771), .B1(n1907), .A0N(sigma15[5]), .A1N(n1938), .Y(
        n1854) );
  XOR2X1 U1800 ( .A(n772), .B(L15_8[5]), .Y(n771) );
  XOR2X1 U1801 ( .A(n773), .B(n774), .Y(n772) );
  OAI2BB2X1 U1802 ( .B0(n35), .B1(n1925), .A0N(sigma5[4]), .A1N(n1929), .Y(
        n1762) );
  XOR2X1 U1803 ( .A(n36), .B(L5_8[4]), .Y(n35) );
  XOR2X1 U1804 ( .A(n37), .B(n38), .Y(n36) );
  OAI2BB2X1 U1805 ( .B0(n971), .B1(n1910), .A0N(sigma12[4]), .A1N(n1942), .Y(
        n1671) );
  XOR2X1 U1806 ( .A(n972), .B(L12_8[4]), .Y(n971) );
  XOR2X1 U1807 ( .A(n973), .B(n974), .Y(n972) );
  OAI2BB2X1 U1808 ( .B0(n2), .B1(n1924), .A0N(sigma5[0]), .A1N(n1934), .Y(
        n1758) );
  XOR2X1 U1809 ( .A(n4), .B(L5_8[0]), .Y(n2) );
  XOR2X1 U1810 ( .A(n5), .B(n6), .Y(n4) );
  OAI2BB2X1 U1811 ( .B0(n43), .B1(n1924), .A0N(sigma5[5]), .A1N(n1931), .Y(
        n1763) );
  XOR2X1 U1812 ( .A(n44), .B(L5_8[5]), .Y(n43) );
  XOR2X1 U1813 ( .A(n45), .B(n46), .Y(n44) );
  OAI2BB2X1 U1814 ( .B0(n251), .B1(n1919), .A0N(sigma3[5]), .A1N(n1946), .Y(
        n1789) );
  XOR2X1 U1815 ( .A(n252), .B(L3_8[5]), .Y(n251) );
  XOR2X1 U1816 ( .A(n253), .B(n254), .Y(n252) );
  OAI2BB2X1 U1817 ( .B0(n347), .B1(n1921), .A0N(sigma2[4]), .A1N(n1942), .Y(
        n1801) );
  XOR2X1 U1818 ( .A(n348), .B(L2_8[4]), .Y(n347) );
  XOR2X1 U1819 ( .A(n349), .B(n350), .Y(n348) );
  OAI2BB2X1 U1820 ( .B0(n667), .B1(n1906), .A0N(sigma14[5]), .A1N(n1936), .Y(
        n1841) );
  XOR2X1 U1821 ( .A(n668), .B(L14_8[5]), .Y(n667) );
  XOR2X1 U1822 ( .A(n669), .B(n670), .Y(n668) );
  OAI2BB2X1 U1823 ( .B0(n1595), .B1(n1918), .A0N(sigma6[4]), .A1N(n1930), .Y(
        n1749) );
  XOR2X1 U1824 ( .A(n1596), .B(L6_8[4]), .Y(n1595) );
  XOR2X1 U1825 ( .A(n1597), .B(n1598), .Y(n1596) );
  OAI2BB2X1 U1826 ( .B0(n1387), .B1(n1915), .A0N(sigma8[4]), .A1N(n1931), .Y(
        n1723) );
  XOR2X1 U1827 ( .A(n1388), .B(L8_8[4]), .Y(n1387) );
  XOR2X1 U1828 ( .A(n1389), .B(n1390), .Y(n1388) );
  OAI2BB2X1 U1829 ( .B0(n723), .B1(n1907), .A0N(sigma14[12]), .A1N(n1937), .Y(
        n1848) );
  XOR2X1 U1830 ( .A(n724), .B(L14_8[12]), .Y(n723) );
  XOR2X1 U1831 ( .A(n725), .B(n726), .Y(n724) );
  OAI2BB2X1 U1832 ( .B0(n1603), .B1(n1918), .A0N(sigma6[5]), .A1N(n1929), .Y(
        n1750) );
  XOR2X1 U1833 ( .A(n1604), .B(L6_8[5]), .Y(n1603) );
  XOR2X1 U1834 ( .A(n1605), .B(n1606), .Y(n1604) );
  OAI2BB2X1 U1835 ( .B0(n243), .B1(n1918), .A0N(sigma3[4]), .A1N(n1946), .Y(
        n1788) );
  XOR2X1 U1836 ( .A(n244), .B(L3_8[4]), .Y(n243) );
  XOR2X1 U1837 ( .A(n245), .B(n246), .Y(n244) );
  OAI2BB2X1 U1838 ( .B0(n1179), .B1(n1912), .A0N(sigma10[4]), .A1N(n1946), .Y(
        n1697) );
  XOR2X1 U1839 ( .A(n1180), .B(L10_8[4]), .Y(n1179) );
  XOR2X1 U1840 ( .A(n1181), .B(n1182), .Y(n1180) );
  OAI2BB2X1 U1841 ( .B0(n659), .B1(n1906), .A0N(sigma14[4]), .A1N(n1936), .Y(
        n1840) );
  XOR2X1 U1842 ( .A(n660), .B(L14_8[4]), .Y(n659) );
  XOR2X1 U1843 ( .A(n661), .B(n662), .Y(n660) );
  OAI2BB2X1 U1844 ( .B0(n1499), .B1(n1916), .A0N(sigma7[5]), .A1N(n1934), .Y(
        n1737) );
  XOR2X1 U1845 ( .A(n1500), .B(L7_8[5]), .Y(n1499) );
  XOR2X1 U1846 ( .A(n1501), .B(n1502), .Y(n1500) );
  OAI2BB2X1 U1847 ( .B0(n355), .B1(n1921), .A0N(sigma2[5]), .A1N(n1942), .Y(
        n1802) );
  XOR2X1 U1848 ( .A(n356), .B(L2_8[5]), .Y(n355) );
  XOR2X1 U1849 ( .A(n357), .B(n358), .Y(n356) );
  OAI2BB2X1 U1850 ( .B0(n451), .B1(n1923), .A0N(sigma1[4]), .A1N(n1938), .Y(
        n1814) );
  XOR2X1 U1851 ( .A(n452), .B(L1_8[4]), .Y(n451) );
  XOR2X1 U1852 ( .A(n453), .B(n454), .Y(n452) );
  OAI2BB2X1 U1853 ( .B0(n939), .B1(n1909), .A0N(sigma12[0]), .A1N(n1941), .Y(
        n1667) );
  XOR2X1 U1854 ( .A(n940), .B(L12_8[0]), .Y(n939) );
  XOR2X1 U1855 ( .A(n941), .B(n942), .Y(n940) );
  OAI2BB2X1 U1856 ( .B0(n1635), .B1(n1918), .A0N(sigma6[9]), .A1N(n1927), .Y(
        n1754) );
  XOR2X1 U1857 ( .A(n1636), .B(L6_8[9]), .Y(n1635) );
  XOR2X1 U1858 ( .A(n1637), .B(n1638), .Y(n1636) );
  OAI2BB2X1 U1859 ( .B0(n1075), .B1(n1911), .A0N(sigma11[4]), .A1N(n1944), .Y(
        n1684) );
  XOR2X1 U1860 ( .A(n1076), .B(L11_8[4]), .Y(n1075) );
  XOR2X1 U1861 ( .A(n1077), .B(n1078), .Y(n1076) );
  OAI2BB2X1 U1862 ( .B0(n627), .B1(n1905), .A0N(sigma14[0]), .A1N(n1935), .Y(
        n1836) );
  XOR2X1 U1863 ( .A(n628), .B(L14_8[0]), .Y(n627) );
  XOR2X1 U1864 ( .A(n629), .B(n630), .Y(n628) );
  OAI2BB2X1 U1865 ( .B0(n915), .B1(n1909), .A0N(sigma13[10]), .A1N(n1941), .Y(
        n1872) );
  XOR2X1 U1866 ( .A(n916), .B(L13_8[10]), .Y(n915) );
  XOR2X1 U1867 ( .A(n917), .B(n918), .Y(n916) );
  XOR2X1 U1868 ( .A(n921), .B(n922), .Y(n917) );
  OAI2BB2X1 U1869 ( .B0(n1043), .B1(n1911), .A0N(sigma11[0]), .A1N(n1943), .Y(
        n1680) );
  XOR2X1 U1870 ( .A(n1044), .B(L11_8[0]), .Y(n1043) );
  XOR2X1 U1871 ( .A(n1045), .B(n1046), .Y(n1044) );
  OAI2BB2X1 U1872 ( .B0(n459), .B1(n1923), .A0N(sigma1[5]), .A1N(n1938), .Y(
        n1815) );
  XOR2X1 U1873 ( .A(n460), .B(L1_8[5]), .Y(n459) );
  XOR2X1 U1874 ( .A(n461), .B(n462), .Y(n460) );
  OAI2BB2X1 U1875 ( .B0(n99), .B1(n1922), .A0N(sigma5[12]), .A1N(n1933), .Y(
        n1770) );
  XOR2X1 U1876 ( .A(n100), .B(L5_8[12]), .Y(n99) );
  XOR2X1 U1877 ( .A(n101), .B(n102), .Y(n100) );
  XOR2X1 U1878 ( .A(n103), .B(n104), .Y(n102) );
  OAI2BB2X1 U1879 ( .B0(n139), .B1(n1921), .A0N(sigma4[4]), .A1N(n1931), .Y(
        n1775) );
  XOR2X1 U1880 ( .A(n140), .B(L4_8[4]), .Y(n139) );
  XOR2X1 U1881 ( .A(n141), .B(n142), .Y(n140) );
  OAI2BB2X1 U1882 ( .B0(n419), .B1(n1922), .A0N(sigma1[0]), .A1N(n1939), .Y(
        n1810) );
  XOR2X1 U1883 ( .A(n420), .B(L1_8[0]), .Y(n419) );
  XOR2X1 U1884 ( .A(n421), .B(n422), .Y(n420) );
  XOR2X1 U1885 ( .A(n425), .B(n426), .Y(n421) );
  XNOR2X1 U1886 ( .A(L2_2[0]), .B(L2_1[0]), .Y(n320) );
  XNOR2X1 U1887 ( .A(L2_2[12]), .B(L2_1[12]), .Y(n416) );
  XNOR2X1 U1888 ( .A(L1_2[11]), .B(L1_1[11]), .Y(n512) );
  XOR2X1 U1889 ( .A(n423), .B(n424), .Y(n422) );
  XNOR2X1 U1890 ( .A(L1_4[0]), .B(L1_3[0]), .Y(n423) );
  XNOR2X1 U1891 ( .A(L1_2[0]), .B(L1_1[0]), .Y(n424) );
  XNOR2X1 U1892 ( .A(L3_2[0]), .B(L3_1[0]), .Y(n216) );
  XNOR2X1 U1893 ( .A(L1_2[2]), .B(L1_1[2]), .Y(n440) );
  XNOR2X1 U1894 ( .A(L1_4[12]), .B(L1_3[12]), .Y(n519) );
  XOR2X1 U1895 ( .A(n521), .B(n522), .Y(n517) );
  XOR2X1 U1896 ( .A(n497), .B(n498), .Y(n493) );
  XNOR2X1 U1897 ( .A(L1_6[9]), .B(L1_5[9]), .Y(n497) );
  XOR2X1 U1898 ( .A(n57), .B(L1_7[9]), .Y(n498) );
  XNOR2X1 U1899 ( .A(L1_2[12]), .B(L1_1[12]), .Y(n520) );
  XNOR2X1 U1900 ( .A(L2_4[12]), .B(L2_3[12]), .Y(n415) );
  OAI2BB2X1 U1901 ( .B0(n595), .B1(n1905), .A0N(sigma16[9]), .A1N(n1935), .Y(
        n1832) );
  XNOR2X1 U1902 ( .A(L5_6[11]), .B(L5_5[11]), .Y(n97) );
  OAI2BB2X1 U1903 ( .B0(n571), .B1(n1905), .A0N(sigma16[6]), .A1N(n1934), .Y(
        n1829) );
  XOR2X1 U1904 ( .A(col0[11]), .B(L13_7[11]), .Y(n930) );
  XOR2X1 U1905 ( .A(n153), .B(L12_7[4]), .Y(n978) );
  XOR2X1 U1906 ( .A(col0[6]), .B(L15_7[6]), .Y(n786) );
  BUFX3 U1907 ( .A(L16_7[2]), .Y(n1903) );
  OAI2BB2X1 U1908 ( .B0(n115), .B1(n1922), .A0N(sigma4[1]), .A1N(n1932), .Y(
        n1772) );
  XNOR2X1 U1909 ( .A(L12_4[4]), .B(L12_3[4]), .Y(n975) );
  XNOR2X1 U1910 ( .A(L15_4[0]), .B(L15_3[0]), .Y(n735) );
  XNOR2X1 U1911 ( .A(L14_4[10]), .B(L14_3[10]), .Y(n711) );
  XOR2X1 U1912 ( .A(n1244), .B(L10_8[12]), .Y(n1243) );
  XOR2X1 U1913 ( .A(n47), .B(L13_7[5]), .Y(n882) );
  XOR2X1 U1914 ( .A(n41), .B(L14_7[12]), .Y(n730) );
  XNOR2XL U1915 ( .A(L4_4[7]), .B(L4_3[7]), .Y(n167) );
  XNOR2X1 U1916 ( .A(L5_4[11]), .B(L5_3[11]), .Y(n95) );
  XNOR2X1 U1917 ( .A(L1_4[9]), .B(L1_3[9]), .Y(n495) );
  XNOR2XL U1918 ( .A(L2_4[0]), .B(L2_3[0]), .Y(n319) );
  XOR2X1 U1919 ( .A(n71), .B(L6_7[2]), .Y(n1586) );
  XNOR2X1 U1920 ( .A(L15_6[7]), .B(L15_5[7]), .Y(n793) );
  XOR2XL U1921 ( .A(col0[3]), .B(L1_7[3]), .Y(n450) );
  XNOR2XL U1922 ( .A(L5_4[2]), .B(L5_3[2]), .Y(n23) );
  XNOR2X1 U1923 ( .A(L3_4[4]), .B(L3_3[4]), .Y(n247) );
  XNOR2XL U1924 ( .A(L5_4[10]), .B(L5_3[10]), .Y(n87) );
  XNOR2XL U1925 ( .A(L6_4[0]), .B(L6_3[0]), .Y(n1567) );
  XOR2X1 U1926 ( .A(n39), .B(L2_7[6]), .Y(n370) );
  XNOR2X1 U1927 ( .A(L16_4[11]), .B(L16_3[11]), .Y(n615) );
  XNOR2X1 U1928 ( .A(L15_4[7]), .B(L15_3[7]), .Y(n791) );
  OAI2BB2X1 U1929 ( .B0(n427), .B1(n1922), .A0N(sigma1[1]), .A1N(n1939), .Y(
        n1811) );
  XOR2XL U1930 ( .A(col0[12]), .B(L1_7[12]), .Y(n522) );
  XOR2X1 U1931 ( .A(n47), .B(L15_7[5]), .Y(n778) );
  XNOR2X1 U1932 ( .A(L11_4[2]), .B(L11_3[2]), .Y(n1063) );
  XNOR2XL U1933 ( .A(L15_6[2]), .B(L15_5[2]), .Y(n753) );
  XNOR2XL U1934 ( .A(L14_6[2]), .B(L14_5[2]), .Y(n649) );
  XOR2XL U1935 ( .A(n116), .B(L4_8[1]), .Y(n115) );
  XNOR2X1 U1936 ( .A(L6_4[7]), .B(L6_3[7]), .Y(n1623) );
  XNOR2X1 U1937 ( .A(L7_4[11]), .B(L7_3[11]), .Y(n1551) );
  OAI2BB2X1 U1938 ( .B0(n1283), .B1(n1914), .A0N(sigma9[4]), .A1N(n1927), .Y(
        n1710) );
  OAI2BB2X1 U1939 ( .B0(n1243), .B1(n1913), .A0N(sigma10[12]), .A1N(n1926), 
        .Y(n1705) );
  XNOR2X1 U1940 ( .A(L2_4[9]), .B(L2_3[9]), .Y(n391) );
  XNOR2X1 U1941 ( .A(L3_4[0]), .B(L3_3[0]), .Y(n215) );
  XNOR2XL U1942 ( .A(L1_6[12]), .B(L1_5[12]), .Y(n521) );
  XNOR2X1 U1943 ( .A(L16_6[3]), .B(L16_5[3]), .Y(n553) );
  XNOR2X1 U1944 ( .A(L15_6[8]), .B(L15_5[8]), .Y(n801) );
  XOR2XL U1945 ( .A(col0[11]), .B(L8_7[11]), .Y(n1450) );
  XOR2XL U1946 ( .A(col0[12]), .B(L13_7[12]), .Y(n938) );
  XOR2X1 U1947 ( .A(n47), .B(L12_7[5]), .Y(n986) );
  XOR2XL U1948 ( .A(n1284), .B(L9_8[4]), .Y(n1283) );
  XNOR2XL U1949 ( .A(L1_4[1]), .B(L1_3[1]), .Y(n431) );
  XOR2XL U1950 ( .A(col0[5]), .B(L1_7[5]), .Y(n466) );
  XOR2XL U1951 ( .A(col0[12]), .B(L2_7[12]), .Y(n418) );
  XNOR2X1 U1952 ( .A(L7_4[12]), .B(L7_3[12]), .Y(n1559) );
  XNOR2X1 U1953 ( .A(L6_4[8]), .B(L6_3[8]), .Y(n1631) );
endmodule


module euclidean_4cells ( deg_Ri, deg_Qi, stop_i, Rin, Qin, Lin, Uin, start, 
        start_cnt, deg_Ro, deg_Qo, stop_o, Rout, Qout, Lout, Uout, st_out, clk, 
        reset );
  input [4:0] deg_Ri;
  input [4:0] deg_Qi;
  input [12:0] Rin;
  input [12:0] Qin;
  input [12:0] Lin;
  input [12:0] Uin;
  output [4:0] deg_Ro;
  output [4:0] deg_Qo;
  output [12:0] Rout;
  output [12:0] Qout;
  output [12:0] Lout;
  output [12:0] Uout;
  input stop_i, start, start_cnt, clk, reset;
  output stop_o, st_out;
  wire   feedback_sel, St_reg, St, SS_reg, START8, SS, Lstop1, LS1, Lstop2,
         LS2, Lstop3, LS3, ST2, out_sel2, START7, START6, START5, START4,
         START3, START2, START1, STOP8, STOP7, STOP6, STOP5, STOP4, STOP3,
         STOP2, STOP1, ST1, N99, N176, N177, N178, N179, N180, N181, N182,
         N183, N184, N185, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n115, n116, n117, n118, n119, n120, n121, n123,
         n124, n125, n126, n127, n128, n129, n131, n132, n133, n134, n135,
         n136, n137, n139, n140, n141, n142, n143, n144, n145, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n163, n164, n165, n166, n167, n168, n169, n171, n172,
         n173, n174, n175, n176, n177, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n319, n320, n321, n322, n323, n324, n325, n327, n329, n330,
         n331, n332, n333, n334, n335, n337, n339, n340, n341, n342, n343,
         n344, n345, n347, n349, n350, n351, n352, n353, n354, n355, n357,
         n359, n360, n361, n362, n363, n364, n365, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n379, n380, n381, n382,
         n383, n384, n385, n387, n389, n390, n391, n392, n393, n394, n395,
         n397, n399, n400, n401, n402, n403, n404, n405, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n645, n648, n651, n654, n663, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n783, n784, n785,
         n786, n787, n788, n789, n791, n792, n793, n794, n795, n796, n797,
         n799, n800, n801, n802, n803, n804, n805, n807, n808, n809, n810,
         n811, n812, n813, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n831, n832, n833, n834,
         n835, n836, n837, n839, n840, n841, n842, n843, n844, n845, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n987, n988, n989, n990, n991,
         n992, n993, n995, n997, n998, n999, n1000, n1001, n1002, n1003, n1005,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1015, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1025, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1055, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1065,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1, n398, n406, n643, n644,
         n646, n647, n649, n650, n652, n653, n655, n656, n657, n658, n659,
         n660, n661, n662, n664, n665, n666, n667, n668, n669, n670, n782,
         n790, n798, n806, n814, n830, n838, n846, n986, n994, n996, n1004,
         n1006, n1014, n1016, n1024, n1026, n1034, n1046, n1054, n1056, n1064,
         n1066, n1074, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432;
  wire   [4:0] dR_reg;
  wire   [4:0] DR8;
  wire   [4:0] dR;
  wire   [4:0] dQ_reg;
  wire   [4:0] DQ8;
  wire   [4:0] dQ;
  wire   [2:0] s_reg;
  wire   [12:0] Rin_reg;
  wire   [12:0] R8;
  wire   [12:0] RR;
  wire   [12:0] Qin_reg;
  wire   [12:0] Q8;
  wire   [12:0] QQ;
  wire   [12:0] Lin_reg;
  wire   [12:0] LLL8;
  wire   [12:0] LL;
  wire   [12:0] Uin_reg;
  wire   [12:0] U8;
  wire   [12:0] UU;
  wire   [4:0] L_dR1;
  wire   [4:0] L_dQ1;
  wire   [12:0] LR1;
  wire   [12:0] LQ1;
  wire   [12:0] LL1;
  wire   [12:0] LU1;
  wire   [2:0] stop1;
  wire   [4:0] L_dR2;
  wire   [4:0] L_dQ2;
  wire   [12:0] LR2;
  wire   [12:0] LQ2;
  wire   [12:0] LL2;
  wire   [12:0] LU2;
  wire   [2:0] stop2;
  wire   [4:0] L_dR3;
  wire   [4:0] L_dQ3;
  wire   [12:0] LR3;
  wire   [12:0] LQ3;
  wire   [12:0] LL3;
  wire   [12:0] LU3;
  wire   [2:0] stop3;
  wire   [12:0] Lout_temp;
  wire   [12:0] out_sel;
  wire   [12:0] L2;
  wire   [12:0] Uout_temp;
  wire   [12:0] U7;
  wire   [12:0] U6;
  wire   [12:0] U5;
  wire   [12:0] U4;
  wire   [12:0] U3;
  wire   [12:0] U2;
  wire   [12:0] U1;
  wire   [12:0] LLL7;
  wire   [12:0] LLL6;
  wire   [12:0] LLL5;
  wire   [12:0] LLL4;
  wire   [12:0] LLL3;
  wire   [12:0] LLL2;
  wire   [12:0] LLL1;
  wire   [12:0] Q7;
  wire   [12:0] Q6;
  wire   [12:0] Q5;
  wire   [12:0] Q4;
  wire   [12:0] Q3;
  wire   [12:0] Q2;
  wire   [12:0] Q1;
  wire   [12:0] R7;
  wire   [12:0] R6;
  wire   [12:0] R5;
  wire   [12:0] R4;
  wire   [12:0] R3;
  wire   [12:0] R2;
  wire   [12:0] R1;
  wire   [4:0] DQ7;
  wire   [4:0] DQ6;
  wire   [4:0] DQ5;
  wire   [4:0] DQ4;
  wire   [4:0] DQ3;
  wire   [4:0] DQ2;
  wire   [4:0] DQ1;
  wire   [4:0] DR7;
  wire   [4:0] DR6;
  wire   [4:0] DR5;
  wire   [4:0] DR4;
  wire   [4:0] DR3;
  wire   [4:0] DR2;
  wire   [4:0] DR1;
  wire   [12:0] L1;
  wire   [9:0] count;
  assign N99 = start_cnt;

  mux_5_2to1_1 mmm1 ( .a(dR_reg), .b(DR8), .sel(n406), .out(dR) );
  mux_5_2to1_0 mmm2 ( .a(dQ_reg), .b(DQ8), .sel(n398), .out(dQ) );
  mux_1_2to1_1 mmm3 ( .a(St_reg), .b(s_reg[2]), .sel(n406), .out(St) );
  mux_13_2to1_3 mmm4 ( .a(Rin_reg), .b(R8), .sel(n398), .out(RR) );
  mux_13_2to1_2 mmm5 ( .a(Qin_reg), .b(Q8), .sel(n398), .out(QQ) );
  mux_13_2to1_1 mmm6 ( .a(Lin_reg), .b(LLL8), .sel(n398), .out(LL) );
  mux_13_2to1_0 mmm7 ( .a(Uin_reg), .b(U8), .sel(feedback_sel), .out(UU) );
  mux_1_2to1_0 mmm8 ( .a(SS_reg), .b(START8), .sel(n406), .out(SS) );
  euclidean_cell_3 cell_1 ( .deg_Ri(dR), .deg_Qi(dQ), .stop_i(St), .Rin(RR), 
        .Qin(QQ), .Lin(LL), .Uin(UU), .start(SS), .start_cnt(n644), .deg_Ro(
        L_dR1), .deg_Qo(L_dQ1), .stop_o(Lstop1), .Rout(LR1), .Qout(LQ1), 
        .Lout(LL1), .Uout(LU1), .st_out(LS1), .clk(clk), .reset(reset) );
  euclidean_cell_2 cell_2 ( .deg_Ri(L_dR1), .deg_Qi(L_dQ1), .stop_i(stop1[2]), 
        .Rin(LR1), .Qin(LQ1), .Lin(LL1), .Uin(LU1), .start(LS1), .start_cnt(
        n1407), .deg_Ro(L_dR2), .deg_Qo(L_dQ2), .stop_o(Lstop2), .Rout(LR2), 
        .Qout(LQ2), .Lout(LL2), .Uout(LU2), .st_out(LS2), .clk(clk), .reset(
        reset) );
  euclidean_cell_1 cell_3 ( .deg_Ri(L_dR2), .deg_Qi(L_dQ2), .stop_i(stop2[2]), 
        .Rin(LR2), .Qin(LQ2), .Lin(LL2), .Uin(LU2), .start(LS2), .start_cnt(
        n643), .deg_Ro(L_dR3), .deg_Qo(L_dQ3), .stop_o(Lstop3), .Rout(LR3), 
        .Qout(LQ3), .Lout(LL3), .Uout(LU3), .st_out(LS3), .clk(clk), .reset(
        reset) );
  euclidean_cell_0 cell_4 ( .deg_Ri(L_dR3), .deg_Qi(L_dQ3), .stop_i(stop3[2]), 
        .Rin(LR3), .Qin(LQ3), .Lin(LL3), .Uin(LU3), .start(LS3), .start_cnt(
        n644), .deg_Ro(deg_Ro), .deg_Qo(deg_Qo), .stop_o(stop_o), .Rout(Rout), 
        .Qout(Qout), .Lout(Lout_temp), .Uout(Uout), .st_out(st_out), .clk(clk), 
        .reset(reset) );
  feedback_ckt_16 F1 ( .Din(Qout), .start(ST2), .Qout(out_sel), .clk(clk), 
        .reset(reset) );
  mux_13_53 m_out ( .a(L2), .b(Uout_temp), .sel(out_sel2), .out(Lout) );
  euclidean_4cells_DW01_inc_0 add_393_S2 ( .A(count), .SUM({N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176}) );
  DFFRHQXL \LLL1_reg[12]  ( .D(n984), .CK(clk), .RN(reset), .Q(LLL1[12]) );
  DFFRHQXL \L1_reg[3]  ( .D(n1410), .CK(clk), .RN(reset), .Q(L1[3]) );
  DFFRHQXL \L1_reg[12]  ( .D(n976), .CK(clk), .RN(reset), .Q(L1[12]) );
  DFFRHQX1 \L1_reg[4]  ( .D(n1412), .CK(clk), .RN(reset), .Q(L1[4]) );
  DFFRHQX1 \R1_reg[5]  ( .D(n1427), .CK(clk), .RN(reset), .Q(R1[5]) );
  DFFRHQXL \L1_reg[5]  ( .D(n1414), .CK(clk), .RN(reset), .Q(L1[5]) );
  DFFRHQXL \L1_reg[7]  ( .D(n1416), .CK(clk), .RN(reset), .Q(L1[7]) );
  DFFRHQX1 \L1_reg[8]  ( .D(n1418), .CK(clk), .RN(reset), .Q(L1[8]) );
  DFFRHQX1 \L1_reg[11]  ( .D(n1424), .CK(clk), .RN(reset), .Q(L1[11]) );
  DFFRHQX1 \R1_reg[3]  ( .D(n1425), .CK(clk), .RN(reset), .Q(R1[3]) );
  DFFRHQX1 \R1_reg[7]  ( .D(n1428), .CK(clk), .RN(reset), .Q(R1[7]) );
  DFFRHQX1 \DR7_reg[4]  ( .D(n675), .CK(clk), .RN(reset), .Q(DR7[4]) );
  DFFRHQX1 \LLL7_reg[0]  ( .D(n1098), .CK(clk), .RN(reset), .Q(LLL7[0]) );
  DFFRHQX1 \LLL7_reg[1]  ( .D(n1088), .CK(clk), .RN(reset), .Q(LLL7[1]) );
  DFFRHQX1 \LLL7_reg[2]  ( .D(n1078), .CK(clk), .RN(reset), .Q(LLL7[2]) );
  DFFRHQX1 \LLL7_reg[3]  ( .D(n1068), .CK(clk), .RN(reset), .Q(LLL7[3]) );
  DFFRHQX1 \LLL7_reg[4]  ( .D(n1058), .CK(clk), .RN(reset), .Q(LLL7[4]) );
  DFFRHQX1 \LLL7_reg[5]  ( .D(n1048), .CK(clk), .RN(reset), .Q(LLL7[5]) );
  DFFRHQX1 \LLL7_reg[6]  ( .D(n1038), .CK(clk), .RN(reset), .Q(LLL7[6]) );
  DFFRHQX1 \LLL7_reg[7]  ( .D(n1028), .CK(clk), .RN(reset), .Q(LLL7[7]) );
  DFFRHQX1 \LLL7_reg[8]  ( .D(n1018), .CK(clk), .RN(reset), .Q(LLL7[8]) );
  DFFRHQX1 \LLL7_reg[9]  ( .D(n1008), .CK(clk), .RN(reset), .Q(LLL7[9]) );
  DFFRHQX1 \LLL7_reg[10]  ( .D(n998), .CK(clk), .RN(reset), .Q(LLL7[10]) );
  DFFRHQX1 \LLL7_reg[11]  ( .D(n988), .CK(clk), .RN(reset), .Q(LLL7[11]) );
  DFFRHQX1 \LLL7_reg[12]  ( .D(n978), .CK(clk), .RN(reset), .Q(LLL7[12]) );
  DFFRHQX1 \Q1_reg[0]  ( .D(n974), .CK(clk), .RN(reset), .Q(Q1[0]) );
  DFFRHQX1 \Q1_reg[1]  ( .D(n966), .CK(clk), .RN(reset), .Q(Q1[1]) );
  DFFRHQX1 \Q1_reg[2]  ( .D(n958), .CK(clk), .RN(reset), .Q(Q1[2]) );
  DFFRHQX1 \Q1_reg[3]  ( .D(n950), .CK(clk), .RN(reset), .Q(Q1[3]) );
  DFFRHQX1 \Q1_reg[4]  ( .D(n942), .CK(clk), .RN(reset), .Q(Q1[4]) );
  DFFRHQX1 \Q1_reg[5]  ( .D(n934), .CK(clk), .RN(reset), .Q(Q1[5]) );
  DFFRHQX1 \Q1_reg[6]  ( .D(n926), .CK(clk), .RN(reset), .Q(Q1[6]) );
  DFFRHQX1 \Q1_reg[7]  ( .D(n918), .CK(clk), .RN(reset), .Q(Q1[7]) );
  DFFRHQX1 \Q1_reg[8]  ( .D(n910), .CK(clk), .RN(reset), .Q(Q1[8]) );
  DFFRHQX1 \Q1_reg[9]  ( .D(n902), .CK(clk), .RN(reset), .Q(Q1[9]) );
  DFFRHQX1 \Q1_reg[10]  ( .D(n894), .CK(clk), .RN(reset), .Q(Q1[10]) );
  DFFRHQX1 \Q1_reg[11]  ( .D(n886), .CK(clk), .RN(reset), .Q(Q1[11]) );
  DFFRHQX1 \Q1_reg[12]  ( .D(n878), .CK(clk), .RN(reset), .Q(Q1[12]) );
  DFFRHQX1 \R1_reg[0]  ( .D(n870), .CK(clk), .RN(reset), .Q(R1[0]) );
  DFFRHQX1 \R1_reg[1]  ( .D(n862), .CK(clk), .RN(reset), .Q(R1[1]) );
  DFFRHQX1 \R1_reg[2]  ( .D(n854), .CK(clk), .RN(reset), .Q(R1[2]) );
  DFFRHQX1 \R1_reg[6]  ( .D(n822), .CK(clk), .RN(reset), .Q(R1[6]) );
  DFFRHQXL \R1_reg[12]  ( .D(n774), .CK(clk), .RN(reset), .Q(R1[12]) );
  DFFRHQX1 \DQ7_reg[0]  ( .D(n747), .CK(clk), .RN(reset), .Q(DQ7[0]) );
  DFFRHQX1 \DQ7_reg[1]  ( .D(n739), .CK(clk), .RN(reset), .Q(DQ7[1]) );
  DFFRHQX1 \DQ7_reg[2]  ( .D(n731), .CK(clk), .RN(reset), .Q(DQ7[2]) );
  DFFRHQX1 \DQ7_reg[3]  ( .D(n723), .CK(clk), .RN(reset), .Q(DQ7[3]) );
  DFFRHQX1 \DQ7_reg[4]  ( .D(n715), .CK(clk), .RN(reset), .Q(DQ7[4]) );
  DFFRHQX1 \DR7_reg[0]  ( .D(n707), .CK(clk), .RN(reset), .Q(DR7[0]) );
  DFFRHQX1 \DR7_reg[1]  ( .D(n699), .CK(clk), .RN(reset), .Q(DR7[1]) );
  DFFRHQX1 \DR7_reg[2]  ( .D(n691), .CK(clk), .RN(reset), .Q(DR7[2]) );
  DFFRHQX1 \DR7_reg[3]  ( .D(n683), .CK(clk), .RN(reset), .Q(DR7[3]) );
  DFFSX1 SS_reg_reg ( .D(n1302), .CK(clk), .SN(reset), .Q(SS_reg), .QN(n672)
         );
  DFFSX1 START8_reg ( .D(n1222), .CK(clk), .SN(reset), .Q(START8), .QN(n663)
         );
  DFFSX1 \stop1_reg[1]  ( .D(n1237), .CK(clk), .SN(reset), .Q(stop1[1]) );
  DFFSX1 \stop2_reg[1]  ( .D(n1234), .CK(clk), .SN(reset), .Q(stop2[1]) );
  DFFSX1 \stop3_reg[1]  ( .D(n1231), .CK(clk), .SN(reset), .Q(stop3[1]) );
  DFFSX1 START7_reg ( .D(n1223), .CK(clk), .SN(reset), .Q(START7) );
  DFFSX1 \s_reg_reg[1]  ( .D(n757), .CK(clk), .SN(reset), .Q(s_reg[1]) );
  DFFSX1 START2_reg ( .D(n1228), .CK(clk), .SN(reset), .Q(START2) );
  DFFSX1 START3_reg ( .D(n1227), .CK(clk), .SN(reset), .Q(START3) );
  DFFSX1 START4_reg ( .D(n1226), .CK(clk), .SN(reset), .Q(START4) );
  DFFSX1 START5_reg ( .D(n1225), .CK(clk), .SN(reset), .Q(START5) );
  DFFSX1 START6_reg ( .D(n1224), .CK(clk), .SN(reset), .Q(START6) );
  DFFSX1 STOP1_reg ( .D(n766), .CK(clk), .SN(reset), .Q(STOP1) );
  DFFSX1 STOP2_reg ( .D(n765), .CK(clk), .SN(reset), .Q(STOP2) );
  DFFSX1 STOP3_reg ( .D(n764), .CK(clk), .SN(reset), .Q(STOP3) );
  DFFSX1 STOP4_reg ( .D(n763), .CK(clk), .SN(reset), .Q(STOP4) );
  DFFSX1 STOP5_reg ( .D(n762), .CK(clk), .SN(reset), .Q(STOP5) );
  DFFSX1 STOP6_reg ( .D(n761), .CK(clk), .SN(reset), .Q(STOP6) );
  DFFSX1 STOP7_reg ( .D(n760), .CK(clk), .SN(reset), .Q(STOP7) );
  DFFSX1 STOP8_reg ( .D(n759), .CK(clk), .SN(reset), .Q(STOP8) );
  DFFSX1 \s_reg_reg[0]  ( .D(n758), .CK(clk), .SN(reset), .Q(s_reg[0]) );
  DFFSX1 \stop1_reg[0]  ( .D(n1238), .CK(clk), .SN(reset), .Q(stop1[0]) );
  DFFSX1 \stop2_reg[0]  ( .D(n1235), .CK(clk), .SN(reset), .Q(stop2[0]) );
  DFFSX1 \stop3_reg[0]  ( .D(n1232), .CK(clk), .SN(reset), .Q(stop3[0]) );
  DFFSX1 START1_reg ( .D(n1229), .CK(clk), .SN(reset), .Q(START1) );
  DFFRHQXL \LLL1_reg[3]  ( .D(n1409), .CK(clk), .RN(reset), .Q(LLL1[3]) );
  DFFRHQX1 \LLL1_reg[4]  ( .D(n1411), .CK(clk), .RN(reset), .Q(LLL1[4]) );
  DFFRHQXL \LLL1_reg[5]  ( .D(n1413), .CK(clk), .RN(reset), .Q(LLL1[5]) );
  DFFRHQXL \LLL1_reg[7]  ( .D(n1415), .CK(clk), .RN(reset), .Q(LLL1[7]) );
  DFFRHQX1 \LLL1_reg[8]  ( .D(n1417), .CK(clk), .RN(reset), .Q(LLL1[8]) );
  DFFRHQX1 \LLL1_reg[11]  ( .D(n1423), .CK(clk), .RN(reset), .Q(LLL1[11]) );
  DFFRHQX1 \Uout_temp_reg[0]  ( .D(n1221), .CK(clk), .RN(reset), .Q(
        Uout_temp[0]) );
  DFFRHQX1 \U8_reg[0]  ( .D(n1213), .CK(clk), .RN(reset), .Q(U8[0]) );
  DFFRHQX1 \Uout_temp_reg[1]  ( .D(n1212), .CK(clk), .RN(reset), .Q(
        Uout_temp[1]) );
  DFFRHQX1 \U8_reg[1]  ( .D(n1204), .CK(clk), .RN(reset), .Q(U8[1]) );
  DFFRHQX1 \Uout_temp_reg[2]  ( .D(n1203), .CK(clk), .RN(reset), .Q(
        Uout_temp[2]) );
  DFFRHQX1 \U8_reg[2]  ( .D(n1195), .CK(clk), .RN(reset), .Q(U8[2]) );
  DFFRHQX1 \Uout_temp_reg[3]  ( .D(n1194), .CK(clk), .RN(reset), .Q(
        Uout_temp[3]) );
  DFFRHQX1 \U8_reg[3]  ( .D(n1186), .CK(clk), .RN(reset), .Q(U8[3]) );
  DFFRHQX1 \Uout_temp_reg[4]  ( .D(n1185), .CK(clk), .RN(reset), .Q(
        Uout_temp[4]) );
  DFFRHQX1 \U8_reg[4]  ( .D(n1177), .CK(clk), .RN(reset), .Q(U8[4]) );
  DFFRHQX1 \Uout_temp_reg[5]  ( .D(n1176), .CK(clk), .RN(reset), .Q(
        Uout_temp[5]) );
  DFFRHQX1 \U8_reg[5]  ( .D(n1168), .CK(clk), .RN(reset), .Q(U8[5]) );
  DFFRHQX1 \Uout_temp_reg[6]  ( .D(n1167), .CK(clk), .RN(reset), .Q(
        Uout_temp[6]) );
  DFFRHQX1 \U8_reg[6]  ( .D(n1159), .CK(clk), .RN(reset), .Q(U8[6]) );
  DFFRHQX1 \Uout_temp_reg[7]  ( .D(n1158), .CK(clk), .RN(reset), .Q(
        Uout_temp[7]) );
  DFFRHQX1 \U8_reg[7]  ( .D(n1150), .CK(clk), .RN(reset), .Q(U8[7]) );
  DFFRHQX1 \Uout_temp_reg[8]  ( .D(n1149), .CK(clk), .RN(reset), .Q(
        Uout_temp[8]) );
  DFFRHQX1 \U8_reg[8]  ( .D(n1141), .CK(clk), .RN(reset), .Q(U8[8]) );
  DFFRHQX1 \Uout_temp_reg[9]  ( .D(n1140), .CK(clk), .RN(reset), .Q(
        Uout_temp[9]) );
  DFFRHQX1 \U8_reg[9]  ( .D(n1132), .CK(clk), .RN(reset), .Q(U8[9]) );
  DFFRHQX1 \Uout_temp_reg[10]  ( .D(n1131), .CK(clk), .RN(reset), .Q(
        Uout_temp[10]) );
  DFFRHQX1 \U8_reg[10]  ( .D(n1123), .CK(clk), .RN(reset), .Q(U8[10]) );
  DFFRHQX1 \Uout_temp_reg[11]  ( .D(n1122), .CK(clk), .RN(reset), .Q(
        Uout_temp[11]) );
  DFFRHQX1 \U8_reg[11]  ( .D(n1114), .CK(clk), .RN(reset), .Q(U8[11]) );
  DFFRHQX1 \Uout_temp_reg[12]  ( .D(n1113), .CK(clk), .RN(reset), .Q(
        Uout_temp[12]) );
  DFFRHQX1 \U8_reg[12]  ( .D(n1105), .CK(clk), .RN(reset), .Q(U8[12]) );
  DFFRHQX1 \LLL8_reg[0]  ( .D(n1097), .CK(clk), .RN(reset), .Q(LLL8[0]) );
  DFFRHQX1 \LLL8_reg[1]  ( .D(n1087), .CK(clk), .RN(reset), .Q(LLL8[1]) );
  DFFRHQX1 \LLL8_reg[2]  ( .D(n1077), .CK(clk), .RN(reset), .Q(LLL8[2]) );
  DFFRHQX1 \LLL8_reg[3]  ( .D(n1067), .CK(clk), .RN(reset), .Q(LLL8[3]) );
  DFFRHQX1 \LLL8_reg[4]  ( .D(n1057), .CK(clk), .RN(reset), .Q(LLL8[4]) );
  DFFRHQX1 \LLL8_reg[5]  ( .D(n1047), .CK(clk), .RN(reset), .Q(LLL8[5]) );
  DFFRHQX1 \LLL8_reg[6]  ( .D(n1037), .CK(clk), .RN(reset), .Q(LLL8[6]) );
  DFFRHQX1 \LLL8_reg[7]  ( .D(n1027), .CK(clk), .RN(reset), .Q(LLL8[7]) );
  DFFRHQX1 \LLL8_reg[8]  ( .D(n1017), .CK(clk), .RN(reset), .Q(LLL8[8]) );
  DFFRHQX1 \LLL8_reg[9]  ( .D(n1007), .CK(clk), .RN(reset), .Q(LLL8[9]) );
  DFFRHQX1 \LLL8_reg[10]  ( .D(n997), .CK(clk), .RN(reset), .Q(LLL8[10]) );
  DFFRHQX1 \LLL8_reg[11]  ( .D(n987), .CK(clk), .RN(reset), .Q(LLL8[11]) );
  DFFRHQX1 \LLL8_reg[12]  ( .D(n977), .CK(clk), .RN(reset), .Q(LLL8[12]) );
  DFFRHQX1 \Q8_reg[0]  ( .D(n967), .CK(clk), .RN(reset), .Q(Q8[0]) );
  DFFRHQX1 \Q8_reg[1]  ( .D(n959), .CK(clk), .RN(reset), .Q(Q8[1]) );
  DFFRHQX1 \Q8_reg[2]  ( .D(n951), .CK(clk), .RN(reset), .Q(Q8[2]) );
  DFFRHQX1 \Q8_reg[3]  ( .D(n943), .CK(clk), .RN(reset), .Q(Q8[3]) );
  DFFRHQX1 \Q8_reg[4]  ( .D(n935), .CK(clk), .RN(reset), .Q(Q8[4]) );
  DFFRHQX1 \Q8_reg[5]  ( .D(n927), .CK(clk), .RN(reset), .Q(Q8[5]) );
  DFFRHQX1 \Q8_reg[6]  ( .D(n919), .CK(clk), .RN(reset), .Q(Q8[6]) );
  DFFRHQX1 \Q8_reg[7]  ( .D(n911), .CK(clk), .RN(reset), .Q(Q8[7]) );
  DFFRHQX1 \Q8_reg[8]  ( .D(n903), .CK(clk), .RN(reset), .Q(Q8[8]) );
  DFFRHQX1 \Q8_reg[9]  ( .D(n895), .CK(clk), .RN(reset), .Q(Q8[9]) );
  DFFRHQX1 \Q8_reg[10]  ( .D(n887), .CK(clk), .RN(reset), .Q(Q8[10]) );
  DFFRHQX1 \Q8_reg[11]  ( .D(n879), .CK(clk), .RN(reset), .Q(Q8[11]) );
  DFFRHQX1 \Q8_reg[12]  ( .D(n871), .CK(clk), .RN(reset), .Q(Q8[12]) );
  DFFRHQX1 \R8_reg[0]  ( .D(n863), .CK(clk), .RN(reset), .Q(R8[0]) );
  DFFRHQX1 \R8_reg[1]  ( .D(n855), .CK(clk), .RN(reset), .Q(R8[1]) );
  DFFRHQX1 \R8_reg[2]  ( .D(n847), .CK(clk), .RN(reset), .Q(R8[2]) );
  DFFRHQX1 \R8_reg[3]  ( .D(n839), .CK(clk), .RN(reset), .Q(R8[3]) );
  DFFRHQX1 \R8_reg[4]  ( .D(n831), .CK(clk), .RN(reset), .Q(R8[4]) );
  DFFRHQX1 \R8_reg[5]  ( .D(n823), .CK(clk), .RN(reset), .Q(R8[5]) );
  DFFRHQX1 \R8_reg[6]  ( .D(n815), .CK(clk), .RN(reset), .Q(R8[6]) );
  DFFRHQX1 \R8_reg[7]  ( .D(n807), .CK(clk), .RN(reset), .Q(R8[7]) );
  DFFRHQX1 \R8_reg[8]  ( .D(n799), .CK(clk), .RN(reset), .Q(R8[8]) );
  DFFRHQX1 \R8_reg[9]  ( .D(n791), .CK(clk), .RN(reset), .Q(R8[9]) );
  DFFRHQX1 \R8_reg[10]  ( .D(n783), .CK(clk), .RN(reset), .Q(R8[10]) );
  DFFRHQX1 \R8_reg[11]  ( .D(n775), .CK(clk), .RN(reset), .Q(R8[11]) );
  DFFRHQX1 \R8_reg[12]  ( .D(n767), .CK(clk), .RN(reset), .Q(R8[12]) );
  DFFRHQX1 \DQ8_reg[0]  ( .D(n746), .CK(clk), .RN(reset), .Q(DQ8[0]) );
  DFFRHQX1 \DQ8_reg[1]  ( .D(n738), .CK(clk), .RN(reset), .Q(DQ8[1]) );
  DFFRHQX1 \DQ8_reg[2]  ( .D(n730), .CK(clk), .RN(reset), .Q(DQ8[2]) );
  DFFRHQX1 \DQ8_reg[4]  ( .D(n714), .CK(clk), .RN(reset), .Q(DQ8[4]) );
  DFFRHQX1 \DR8_reg[0]  ( .D(n706), .CK(clk), .RN(reset), .Q(DR8[0]) );
  DFFRHQX1 \DR8_reg[1]  ( .D(n698), .CK(clk), .RN(reset), .Q(DR8[1]) );
  DFFRHQX1 \DR8_reg[2]  ( .D(n690), .CK(clk), .RN(reset), .Q(DR8[2]) );
  DFFRHQX1 \DR8_reg[3]  ( .D(n682), .CK(clk), .RN(reset), .Q(DR8[3]) );
  DFFRHQX1 \DR8_reg[4]  ( .D(n674), .CK(clk), .RN(reset), .Q(DR8[4]) );
  DFFRHQX1 \LLL1_reg[0]  ( .D(n1104), .CK(clk), .RN(reset), .Q(LLL1[0]) );
  DFFRHQX1 \LLL1_reg[1]  ( .D(n1094), .CK(clk), .RN(reset), .Q(LLL1[1]) );
  DFFRHQX1 \LLL1_reg[2]  ( .D(n1084), .CK(clk), .RN(reset), .Q(LLL1[2]) );
  DFFRHQX1 \LLL1_reg[6]  ( .D(n1044), .CK(clk), .RN(reset), .Q(LLL1[6]) );
  DFFRHQX1 \Lin_reg_reg[12]  ( .D(n1275), .CK(clk), .RN(reset), .Q(Lin_reg[12]) );
  DFFRHQX1 \Lin_reg_reg[11]  ( .D(n1274), .CK(clk), .RN(reset), .Q(Lin_reg[11]) );
  DFFRHQX1 \Lin_reg_reg[10]  ( .D(n1273), .CK(clk), .RN(reset), .Q(Lin_reg[10]) );
  DFFRHQX1 \Lin_reg_reg[8]  ( .D(n1271), .CK(clk), .RN(reset), .Q(Lin_reg[8])
         );
  DFFRHQX1 \Lin_reg_reg[7]  ( .D(n1270), .CK(clk), .RN(reset), .Q(Lin_reg[7])
         );
  DFFRHQX1 \Lin_reg_reg[6]  ( .D(n1269), .CK(clk), .RN(reset), .Q(Lin_reg[6])
         );
  DFFRHQX1 \Lin_reg_reg[5]  ( .D(n1268), .CK(clk), .RN(reset), .Q(Lin_reg[5])
         );
  DFFRHQX1 \Lin_reg_reg[4]  ( .D(n1267), .CK(clk), .RN(reset), .Q(Lin_reg[4])
         );
  DFFRHQX1 \Lin_reg_reg[3]  ( .D(n1266), .CK(clk), .RN(reset), .Q(Lin_reg[3])
         );
  DFFRHQX1 \Lin_reg_reg[2]  ( .D(n1265), .CK(clk), .RN(reset), .Q(Lin_reg[2])
         );
  DFFRHQX1 \Lin_reg_reg[1]  ( .D(n1264), .CK(clk), .RN(reset), .Q(Lin_reg[1])
         );
  DFFRHQX1 \Lin_reg_reg[0]  ( .D(n1263), .CK(clk), .RN(reset), .Q(Lin_reg[0])
         );
  DFFRHQX1 \L2_reg[0]  ( .D(n1095), .CK(clk), .RN(reset), .Q(L2[0]) );
  DFFRHQX1 \L2_reg[1]  ( .D(n1085), .CK(clk), .RN(reset), .Q(L2[1]) );
  DFFRHQX1 \L2_reg[2]  ( .D(n1075), .CK(clk), .RN(reset), .Q(L2[2]) );
  DFFRHQX1 \L2_reg[3]  ( .D(n1065), .CK(clk), .RN(reset), .Q(L2[3]) );
  DFFRHQX1 \L2_reg[4]  ( .D(n1055), .CK(clk), .RN(reset), .Q(L2[4]) );
  DFFRHQX1 \L2_reg[5]  ( .D(n1045), .CK(clk), .RN(reset), .Q(L2[5]) );
  DFFRHQX1 \L2_reg[6]  ( .D(n1035), .CK(clk), .RN(reset), .Q(L2[6]) );
  DFFRHQX1 \L2_reg[7]  ( .D(n1025), .CK(clk), .RN(reset), .Q(L2[7]) );
  DFFRHQX1 \L2_reg[8]  ( .D(n1015), .CK(clk), .RN(reset), .Q(L2[8]) );
  DFFRHQX1 \L2_reg[10]  ( .D(n995), .CK(clk), .RN(reset), .Q(L2[10]) );
  DFFRHQX1 \L2_reg[11]  ( .D(n985), .CK(clk), .RN(reset), .Q(L2[11]) );
  DFFRHQX1 \L2_reg[12]  ( .D(n975), .CK(clk), .RN(reset), .Q(L2[12]) );
  DFFRHQX1 \dR_reg_reg[3]  ( .D(n1312), .CK(clk), .RN(reset), .Q(dR_reg[3]) );
  DFFRHQX1 \dR_reg_reg[2]  ( .D(n1311), .CK(clk), .RN(reset), .Q(dR_reg[2]) );
  DFFRHQX1 \dR_reg_reg[1]  ( .D(n1310), .CK(clk), .RN(reset), .Q(dR_reg[1]) );
  DFFRHQX1 \dR_reg_reg[0]  ( .D(n1309), .CK(clk), .RN(reset), .Q(dR_reg[0]) );
  DFFRHQX1 \dQ_reg_reg[2]  ( .D(n1306), .CK(clk), .RN(reset), .Q(dQ_reg[2]) );
  DFFRHQX1 \dQ_reg_reg[1]  ( .D(n1305), .CK(clk), .RN(reset), .Q(dQ_reg[1]) );
  DFFRHQX1 \dQ_reg_reg[0]  ( .D(n1304), .CK(clk), .RN(reset), .Q(dQ_reg[0]) );
  DFFRHQX1 \Rin_reg_reg[12]  ( .D(n1301), .CK(clk), .RN(reset), .Q(Rin_reg[12]) );
  DFFRHQX1 \Rin_reg_reg[11]  ( .D(n1300), .CK(clk), .RN(reset), .Q(Rin_reg[11]) );
  DFFRHQX1 \Rin_reg_reg[10]  ( .D(n1299), .CK(clk), .RN(reset), .Q(Rin_reg[10]) );
  DFFRHQX1 \Rin_reg_reg[8]  ( .D(n1297), .CK(clk), .RN(reset), .Q(Rin_reg[8])
         );
  DFFRHQX1 \Rin_reg_reg[7]  ( .D(n1296), .CK(clk), .RN(reset), .Q(Rin_reg[7])
         );
  DFFRHQX1 \Rin_reg_reg[6]  ( .D(n1295), .CK(clk), .RN(reset), .Q(Rin_reg[6])
         );
  DFFRHQX1 \Rin_reg_reg[5]  ( .D(n1294), .CK(clk), .RN(reset), .Q(Rin_reg[5])
         );
  DFFRHQX1 \Rin_reg_reg[4]  ( .D(n1293), .CK(clk), .RN(reset), .Q(Rin_reg[4])
         );
  DFFRHQX1 \Rin_reg_reg[3]  ( .D(n1292), .CK(clk), .RN(reset), .Q(Rin_reg[3])
         );
  DFFRHQX1 \Rin_reg_reg[2]  ( .D(n1291), .CK(clk), .RN(reset), .Q(Rin_reg[2])
         );
  DFFRHQX1 \Rin_reg_reg[1]  ( .D(n1290), .CK(clk), .RN(reset), .Q(Rin_reg[1])
         );
  DFFRHQX1 \Rin_reg_reg[0]  ( .D(n1289), .CK(clk), .RN(reset), .Q(Rin_reg[0])
         );
  DFFRHQX1 \Qin_reg_reg[12]  ( .D(n1288), .CK(clk), .RN(reset), .Q(Qin_reg[12]) );
  DFFRHQX1 \Qin_reg_reg[11]  ( .D(n1287), .CK(clk), .RN(reset), .Q(Qin_reg[11]) );
  DFFRHQX1 \Qin_reg_reg[10]  ( .D(n1286), .CK(clk), .RN(reset), .Q(Qin_reg[10]) );
  DFFRHQX1 \Qin_reg_reg[8]  ( .D(n1284), .CK(clk), .RN(reset), .Q(Qin_reg[8])
         );
  DFFRHQX1 \Qin_reg_reg[7]  ( .D(n1283), .CK(clk), .RN(reset), .Q(Qin_reg[7])
         );
  DFFRHQX1 \Qin_reg_reg[6]  ( .D(n1282), .CK(clk), .RN(reset), .Q(Qin_reg[6])
         );
  DFFRHQX1 \Qin_reg_reg[5]  ( .D(n1281), .CK(clk), .RN(reset), .Q(Qin_reg[5])
         );
  DFFRHQX1 \Qin_reg_reg[4]  ( .D(n1280), .CK(clk), .RN(reset), .Q(Qin_reg[4])
         );
  DFFRHQX1 \Qin_reg_reg[3]  ( .D(n1279), .CK(clk), .RN(reset), .Q(Qin_reg[3])
         );
  DFFRHQX1 \Qin_reg_reg[2]  ( .D(n1278), .CK(clk), .RN(reset), .Q(Qin_reg[2])
         );
  DFFRHQX1 \Qin_reg_reg[1]  ( .D(n1277), .CK(clk), .RN(reset), .Q(Qin_reg[1])
         );
  DFFRHQX1 \Qin_reg_reg[0]  ( .D(n1276), .CK(clk), .RN(reset), .Q(Qin_reg[0])
         );
  DFFRHQX1 \Uin_reg_reg[12]  ( .D(n1262), .CK(clk), .RN(reset), .Q(Uin_reg[12]) );
  DFFRHQX1 \Uin_reg_reg[11]  ( .D(n1261), .CK(clk), .RN(reset), .Q(Uin_reg[11]) );
  DFFRHQX1 \Uin_reg_reg[10]  ( .D(n1260), .CK(clk), .RN(reset), .Q(Uin_reg[10]) );
  DFFRHQX1 \Uin_reg_reg[8]  ( .D(n1258), .CK(clk), .RN(reset), .Q(Uin_reg[8])
         );
  DFFRHQX1 \Uin_reg_reg[7]  ( .D(n1257), .CK(clk), .RN(reset), .Q(Uin_reg[7])
         );
  DFFRHQX1 \Uin_reg_reg[6]  ( .D(n1256), .CK(clk), .RN(reset), .Q(Uin_reg[6])
         );
  DFFRHQX1 \Uin_reg_reg[5]  ( .D(n1255), .CK(clk), .RN(reset), .Q(Uin_reg[5])
         );
  DFFRHQX1 \Uin_reg_reg[4]  ( .D(n1254), .CK(clk), .RN(reset), .Q(Uin_reg[4])
         );
  DFFRHQX1 \Uin_reg_reg[3]  ( .D(n1253), .CK(clk), .RN(reset), .Q(Uin_reg[3])
         );
  DFFRHQX1 \Uin_reg_reg[2]  ( .D(n1252), .CK(clk), .RN(reset), .Q(Uin_reg[2])
         );
  DFFRHQX1 \Uin_reg_reg[1]  ( .D(n1251), .CK(clk), .RN(reset), .Q(Uin_reg[1])
         );
  DFFRHQX1 \Uin_reg_reg[0]  ( .D(n1250), .CK(clk), .RN(reset), .Q(Uin_reg[0])
         );
  DFFRHQX1 \Lin_reg_reg[9]  ( .D(n1272), .CK(clk), .RN(reset), .Q(Lin_reg[9])
         );
  DFFRHQX1 \L2_reg[9]  ( .D(n1005), .CK(clk), .RN(reset), .Q(L2[9]) );
  DFFRHQX1 \U1_reg[0]  ( .D(n1220), .CK(clk), .RN(reset), .Q(U1[0]) );
  DFFRHQX1 \U2_reg[0]  ( .D(n1219), .CK(clk), .RN(reset), .Q(U2[0]) );
  DFFRHQX1 \U3_reg[0]  ( .D(n1218), .CK(clk), .RN(reset), .Q(U3[0]) );
  DFFRHQX1 \U4_reg[0]  ( .D(n1217), .CK(clk), .RN(reset), .Q(U4[0]) );
  DFFRHQX1 \U5_reg[0]  ( .D(n1216), .CK(clk), .RN(reset), .Q(U5[0]) );
  DFFRHQX1 \U6_reg[0]  ( .D(n1215), .CK(clk), .RN(reset), .Q(U6[0]) );
  DFFRHQX1 \U7_reg[0]  ( .D(n1214), .CK(clk), .RN(reset), .Q(U7[0]) );
  DFFRHQX1 \U1_reg[1]  ( .D(n1211), .CK(clk), .RN(reset), .Q(U1[1]) );
  DFFRHQX1 \U2_reg[1]  ( .D(n1210), .CK(clk), .RN(reset), .Q(U2[1]) );
  DFFRHQX1 \U3_reg[1]  ( .D(n1209), .CK(clk), .RN(reset), .Q(U3[1]) );
  DFFRHQX1 \U4_reg[1]  ( .D(n1208), .CK(clk), .RN(reset), .Q(U4[1]) );
  DFFRHQX1 \U5_reg[1]  ( .D(n1207), .CK(clk), .RN(reset), .Q(U5[1]) );
  DFFRHQX1 \U6_reg[1]  ( .D(n1206), .CK(clk), .RN(reset), .Q(U6[1]) );
  DFFRHQX1 \U7_reg[1]  ( .D(n1205), .CK(clk), .RN(reset), .Q(U7[1]) );
  DFFRHQX1 \U1_reg[2]  ( .D(n1202), .CK(clk), .RN(reset), .Q(U1[2]) );
  DFFRHQX1 \U2_reg[2]  ( .D(n1201), .CK(clk), .RN(reset), .Q(U2[2]) );
  DFFRHQX1 \U3_reg[2]  ( .D(n1200), .CK(clk), .RN(reset), .Q(U3[2]) );
  DFFRHQX1 \U4_reg[2]  ( .D(n1199), .CK(clk), .RN(reset), .Q(U4[2]) );
  DFFRHQX1 \U5_reg[2]  ( .D(n1198), .CK(clk), .RN(reset), .Q(U5[2]) );
  DFFRHQX1 \U6_reg[2]  ( .D(n1197), .CK(clk), .RN(reset), .Q(U6[2]) );
  DFFRHQX1 \U7_reg[2]  ( .D(n1196), .CK(clk), .RN(reset), .Q(U7[2]) );
  DFFRHQX1 \U1_reg[3]  ( .D(n1193), .CK(clk), .RN(reset), .Q(U1[3]) );
  DFFRHQX1 \U2_reg[3]  ( .D(n1192), .CK(clk), .RN(reset), .Q(U2[3]) );
  DFFRHQX1 \U3_reg[3]  ( .D(n1191), .CK(clk), .RN(reset), .Q(U3[3]) );
  DFFRHQX1 \U4_reg[3]  ( .D(n1190), .CK(clk), .RN(reset), .Q(U4[3]) );
  DFFRHQX1 \U5_reg[3]  ( .D(n1189), .CK(clk), .RN(reset), .Q(U5[3]) );
  DFFRHQX1 \U6_reg[3]  ( .D(n1188), .CK(clk), .RN(reset), .Q(U6[3]) );
  DFFRHQX1 \U7_reg[3]  ( .D(n1187), .CK(clk), .RN(reset), .Q(U7[3]) );
  DFFRHQX1 \U1_reg[4]  ( .D(n1184), .CK(clk), .RN(reset), .Q(U1[4]) );
  DFFRHQX1 \U2_reg[4]  ( .D(n1183), .CK(clk), .RN(reset), .Q(U2[4]) );
  DFFRHQX1 \U3_reg[4]  ( .D(n1182), .CK(clk), .RN(reset), .Q(U3[4]) );
  DFFRHQX1 \U4_reg[4]  ( .D(n1181), .CK(clk), .RN(reset), .Q(U4[4]) );
  DFFRHQX1 \U5_reg[4]  ( .D(n1180), .CK(clk), .RN(reset), .Q(U5[4]) );
  DFFRHQX1 \U6_reg[4]  ( .D(n1179), .CK(clk), .RN(reset), .Q(U6[4]) );
  DFFRHQX1 \U7_reg[4]  ( .D(n1178), .CK(clk), .RN(reset), .Q(U7[4]) );
  DFFRHQX1 \U1_reg[5]  ( .D(n1175), .CK(clk), .RN(reset), .Q(U1[5]) );
  DFFRHQX1 \U2_reg[5]  ( .D(n1174), .CK(clk), .RN(reset), .Q(U2[5]) );
  DFFRHQX1 \U3_reg[5]  ( .D(n1173), .CK(clk), .RN(reset), .Q(U3[5]) );
  DFFRHQX1 \U4_reg[5]  ( .D(n1172), .CK(clk), .RN(reset), .Q(U4[5]) );
  DFFRHQX1 \U5_reg[5]  ( .D(n1171), .CK(clk), .RN(reset), .Q(U5[5]) );
  DFFRHQX1 \U6_reg[5]  ( .D(n1170), .CK(clk), .RN(reset), .Q(U6[5]) );
  DFFRHQX1 \U7_reg[5]  ( .D(n1169), .CK(clk), .RN(reset), .Q(U7[5]) );
  DFFRHQX1 \U1_reg[6]  ( .D(n1166), .CK(clk), .RN(reset), .Q(U1[6]) );
  DFFRHQX1 \U2_reg[6]  ( .D(n1165), .CK(clk), .RN(reset), .Q(U2[6]) );
  DFFRHQX1 \U3_reg[6]  ( .D(n1164), .CK(clk), .RN(reset), .Q(U3[6]) );
  DFFRHQX1 \U4_reg[6]  ( .D(n1163), .CK(clk), .RN(reset), .Q(U4[6]) );
  DFFRHQX1 \U5_reg[6]  ( .D(n1162), .CK(clk), .RN(reset), .Q(U5[6]) );
  DFFRHQX1 \U6_reg[6]  ( .D(n1161), .CK(clk), .RN(reset), .Q(U6[6]) );
  DFFRHQX1 \U7_reg[6]  ( .D(n1160), .CK(clk), .RN(reset), .Q(U7[6]) );
  DFFRHQX1 \U1_reg[7]  ( .D(n1157), .CK(clk), .RN(reset), .Q(U1[7]) );
  DFFRHQX1 \U2_reg[7]  ( .D(n1156), .CK(clk), .RN(reset), .Q(U2[7]) );
  DFFRHQX1 \U3_reg[7]  ( .D(n1155), .CK(clk), .RN(reset), .Q(U3[7]) );
  DFFRHQX1 \U4_reg[7]  ( .D(n1154), .CK(clk), .RN(reset), .Q(U4[7]) );
  DFFRHQX1 \U5_reg[7]  ( .D(n1153), .CK(clk), .RN(reset), .Q(U5[7]) );
  DFFRHQX1 \U6_reg[7]  ( .D(n1152), .CK(clk), .RN(reset), .Q(U6[7]) );
  DFFRHQX1 \U7_reg[7]  ( .D(n1151), .CK(clk), .RN(reset), .Q(U7[7]) );
  DFFRHQX1 \U1_reg[8]  ( .D(n1148), .CK(clk), .RN(reset), .Q(U1[8]) );
  DFFRHQX1 \U2_reg[8]  ( .D(n1147), .CK(clk), .RN(reset), .Q(U2[8]) );
  DFFRHQX1 \U3_reg[8]  ( .D(n1146), .CK(clk), .RN(reset), .Q(U3[8]) );
  DFFRHQX1 \U4_reg[8]  ( .D(n1145), .CK(clk), .RN(reset), .Q(U4[8]) );
  DFFRHQX1 \U5_reg[8]  ( .D(n1144), .CK(clk), .RN(reset), .Q(U5[8]) );
  DFFRHQX1 \U6_reg[8]  ( .D(n1143), .CK(clk), .RN(reset), .Q(U6[8]) );
  DFFRHQX1 \U7_reg[8]  ( .D(n1142), .CK(clk), .RN(reset), .Q(U7[8]) );
  DFFRHQX1 \U1_reg[9]  ( .D(n1139), .CK(clk), .RN(reset), .Q(U1[9]) );
  DFFRHQX1 \U2_reg[9]  ( .D(n1138), .CK(clk), .RN(reset), .Q(U2[9]) );
  DFFRHQX1 \U3_reg[9]  ( .D(n1137), .CK(clk), .RN(reset), .Q(U3[9]) );
  DFFRHQX1 \U4_reg[9]  ( .D(n1136), .CK(clk), .RN(reset), .Q(U4[9]) );
  DFFRHQX1 \U5_reg[9]  ( .D(n1135), .CK(clk), .RN(reset), .Q(U5[9]) );
  DFFRHQX1 \U6_reg[9]  ( .D(n1134), .CK(clk), .RN(reset), .Q(U6[9]) );
  DFFRHQX1 \U7_reg[9]  ( .D(n1133), .CK(clk), .RN(reset), .Q(U7[9]) );
  DFFRHQX1 \U1_reg[10]  ( .D(n1130), .CK(clk), .RN(reset), .Q(U1[10]) );
  DFFRHQX1 \U2_reg[10]  ( .D(n1129), .CK(clk), .RN(reset), .Q(U2[10]) );
  DFFRHQX1 \U3_reg[10]  ( .D(n1128), .CK(clk), .RN(reset), .Q(U3[10]) );
  DFFRHQX1 \U4_reg[10]  ( .D(n1127), .CK(clk), .RN(reset), .Q(U4[10]) );
  DFFRHQX1 \U5_reg[10]  ( .D(n1126), .CK(clk), .RN(reset), .Q(U5[10]) );
  DFFRHQX1 \U6_reg[10]  ( .D(n1125), .CK(clk), .RN(reset), .Q(U6[10]) );
  DFFRHQX1 \U7_reg[10]  ( .D(n1124), .CK(clk), .RN(reset), .Q(U7[10]) );
  DFFRHQX1 \U1_reg[11]  ( .D(n1121), .CK(clk), .RN(reset), .Q(U1[11]) );
  DFFRHQX1 \U2_reg[11]  ( .D(n1120), .CK(clk), .RN(reset), .Q(U2[11]) );
  DFFRHQX1 \U3_reg[11]  ( .D(n1119), .CK(clk), .RN(reset), .Q(U3[11]) );
  DFFRHQX1 \U4_reg[11]  ( .D(n1118), .CK(clk), .RN(reset), .Q(U4[11]) );
  DFFRHQX1 \U5_reg[11]  ( .D(n1117), .CK(clk), .RN(reset), .Q(U5[11]) );
  DFFRHQX1 \U6_reg[11]  ( .D(n1116), .CK(clk), .RN(reset), .Q(U6[11]) );
  DFFRHQX1 \U7_reg[11]  ( .D(n1115), .CK(clk), .RN(reset), .Q(U7[11]) );
  DFFRHQX1 \U1_reg[12]  ( .D(n1112), .CK(clk), .RN(reset), .Q(U1[12]) );
  DFFRHQX1 \U2_reg[12]  ( .D(n1111), .CK(clk), .RN(reset), .Q(U2[12]) );
  DFFRHQX1 \U3_reg[12]  ( .D(n1110), .CK(clk), .RN(reset), .Q(U3[12]) );
  DFFRHQX1 \U4_reg[12]  ( .D(n1109), .CK(clk), .RN(reset), .Q(U4[12]) );
  DFFRHQX1 \U5_reg[12]  ( .D(n1108), .CK(clk), .RN(reset), .Q(U5[12]) );
  DFFRHQX1 \U6_reg[12]  ( .D(n1107), .CK(clk), .RN(reset), .Q(U6[12]) );
  DFFRHQX1 \U7_reg[12]  ( .D(n1106), .CK(clk), .RN(reset), .Q(U7[12]) );
  DFFRHQX1 \LLL2_reg[0]  ( .D(n1103), .CK(clk), .RN(reset), .Q(LLL2[0]) );
  DFFRHQX1 \LLL3_reg[0]  ( .D(n1102), .CK(clk), .RN(reset), .Q(LLL3[0]) );
  DFFRHQX1 \LLL4_reg[0]  ( .D(n1101), .CK(clk), .RN(reset), .Q(LLL4[0]) );
  DFFRHQX1 \LLL5_reg[0]  ( .D(n1100), .CK(clk), .RN(reset), .Q(LLL5[0]) );
  DFFRHQX1 \LLL6_reg[0]  ( .D(n1099), .CK(clk), .RN(reset), .Q(LLL6[0]) );
  DFFRHQX1 \L1_reg[0]  ( .D(n1096), .CK(clk), .RN(reset), .Q(L1[0]) );
  DFFRHQX1 \LLL2_reg[1]  ( .D(n1093), .CK(clk), .RN(reset), .Q(LLL2[1]) );
  DFFRHQX1 \LLL3_reg[1]  ( .D(n1092), .CK(clk), .RN(reset), .Q(LLL3[1]) );
  DFFRHQX1 \LLL4_reg[1]  ( .D(n1091), .CK(clk), .RN(reset), .Q(LLL4[1]) );
  DFFRHQX1 \LLL5_reg[1]  ( .D(n1090), .CK(clk), .RN(reset), .Q(LLL5[1]) );
  DFFRHQX1 \LLL6_reg[1]  ( .D(n1089), .CK(clk), .RN(reset), .Q(LLL6[1]) );
  DFFRHQX1 \L1_reg[1]  ( .D(n1086), .CK(clk), .RN(reset), .Q(L1[1]) );
  DFFRHQX1 \LLL2_reg[2]  ( .D(n1083), .CK(clk), .RN(reset), .Q(LLL2[2]) );
  DFFRHQX1 \LLL3_reg[2]  ( .D(n1082), .CK(clk), .RN(reset), .Q(LLL3[2]) );
  DFFRHQX1 \LLL4_reg[2]  ( .D(n1081), .CK(clk), .RN(reset), .Q(LLL4[2]) );
  DFFRHQX1 \LLL5_reg[2]  ( .D(n1080), .CK(clk), .RN(reset), .Q(LLL5[2]) );
  DFFRHQX1 \LLL6_reg[2]  ( .D(n1079), .CK(clk), .RN(reset), .Q(LLL6[2]) );
  DFFRHQX1 \L1_reg[2]  ( .D(n1076), .CK(clk), .RN(reset), .Q(L1[2]) );
  DFFRHQX1 \LLL2_reg[3]  ( .D(n1073), .CK(clk), .RN(reset), .Q(LLL2[3]) );
  DFFRHQX1 \LLL3_reg[3]  ( .D(n1072), .CK(clk), .RN(reset), .Q(LLL3[3]) );
  DFFRHQX1 \LLL4_reg[3]  ( .D(n1071), .CK(clk), .RN(reset), .Q(LLL4[3]) );
  DFFRHQX1 \LLL5_reg[3]  ( .D(n1070), .CK(clk), .RN(reset), .Q(LLL5[3]) );
  DFFRHQX1 \LLL6_reg[3]  ( .D(n1069), .CK(clk), .RN(reset), .Q(LLL6[3]) );
  DFFRHQX1 \LLL2_reg[4]  ( .D(n1063), .CK(clk), .RN(reset), .Q(LLL2[4]) );
  DFFRHQX1 \LLL3_reg[4]  ( .D(n1062), .CK(clk), .RN(reset), .Q(LLL3[4]) );
  DFFRHQX1 \LLL4_reg[4]  ( .D(n1061), .CK(clk), .RN(reset), .Q(LLL4[4]) );
  DFFRHQX1 \LLL5_reg[4]  ( .D(n1060), .CK(clk), .RN(reset), .Q(LLL5[4]) );
  DFFRHQX1 \LLL6_reg[4]  ( .D(n1059), .CK(clk), .RN(reset), .Q(LLL6[4]) );
  DFFRHQX1 \LLL2_reg[5]  ( .D(n1053), .CK(clk), .RN(reset), .Q(LLL2[5]) );
  DFFRHQX1 \LLL3_reg[5]  ( .D(n1052), .CK(clk), .RN(reset), .Q(LLL3[5]) );
  DFFRHQX1 \LLL4_reg[5]  ( .D(n1051), .CK(clk), .RN(reset), .Q(LLL4[5]) );
  DFFRHQX1 \LLL5_reg[5]  ( .D(n1050), .CK(clk), .RN(reset), .Q(LLL5[5]) );
  DFFRHQX1 \LLL6_reg[5]  ( .D(n1049), .CK(clk), .RN(reset), .Q(LLL6[5]) );
  DFFRHQX1 \LLL2_reg[6]  ( .D(n1043), .CK(clk), .RN(reset), .Q(LLL2[6]) );
  DFFRHQX1 \LLL3_reg[6]  ( .D(n1042), .CK(clk), .RN(reset), .Q(LLL3[6]) );
  DFFRHQX1 \LLL4_reg[6]  ( .D(n1041), .CK(clk), .RN(reset), .Q(LLL4[6]) );
  DFFRHQX1 \LLL5_reg[6]  ( .D(n1040), .CK(clk), .RN(reset), .Q(LLL5[6]) );
  DFFRHQX1 \LLL6_reg[6]  ( .D(n1039), .CK(clk), .RN(reset), .Q(LLL6[6]) );
  DFFRHQX1 \L1_reg[6]  ( .D(n1036), .CK(clk), .RN(reset), .Q(L1[6]) );
  DFFRHQX1 \LLL2_reg[7]  ( .D(n1033), .CK(clk), .RN(reset), .Q(LLL2[7]) );
  DFFRHQX1 \LLL3_reg[7]  ( .D(n1032), .CK(clk), .RN(reset), .Q(LLL3[7]) );
  DFFRHQX1 \LLL4_reg[7]  ( .D(n1031), .CK(clk), .RN(reset), .Q(LLL4[7]) );
  DFFRHQX1 \LLL5_reg[7]  ( .D(n1030), .CK(clk), .RN(reset), .Q(LLL5[7]) );
  DFFRHQX1 \LLL6_reg[7]  ( .D(n1029), .CK(clk), .RN(reset), .Q(LLL6[7]) );
  DFFRHQX1 \LLL2_reg[8]  ( .D(n1023), .CK(clk), .RN(reset), .Q(LLL2[8]) );
  DFFRHQX1 \LLL3_reg[8]  ( .D(n1022), .CK(clk), .RN(reset), .Q(LLL3[8]) );
  DFFRHQX1 \LLL4_reg[8]  ( .D(n1021), .CK(clk), .RN(reset), .Q(LLL4[8]) );
  DFFRHQX1 \LLL5_reg[8]  ( .D(n1020), .CK(clk), .RN(reset), .Q(LLL5[8]) );
  DFFRHQX1 \LLL6_reg[8]  ( .D(n1019), .CK(clk), .RN(reset), .Q(LLL6[8]) );
  DFFRHQX1 \LLL2_reg[9]  ( .D(n1013), .CK(clk), .RN(reset), .Q(LLL2[9]) );
  DFFRHQX1 \LLL3_reg[9]  ( .D(n1012), .CK(clk), .RN(reset), .Q(LLL3[9]) );
  DFFRHQX1 \LLL4_reg[9]  ( .D(n1011), .CK(clk), .RN(reset), .Q(LLL4[9]) );
  DFFRHQX1 \LLL5_reg[9]  ( .D(n1010), .CK(clk), .RN(reset), .Q(LLL5[9]) );
  DFFRHQX1 \LLL6_reg[9]  ( .D(n1009), .CK(clk), .RN(reset), .Q(LLL6[9]) );
  DFFRHQX1 \LLL2_reg[10]  ( .D(n1003), .CK(clk), .RN(reset), .Q(LLL2[10]) );
  DFFRHQX1 \LLL3_reg[10]  ( .D(n1002), .CK(clk), .RN(reset), .Q(LLL3[10]) );
  DFFRHQX1 \LLL4_reg[10]  ( .D(n1001), .CK(clk), .RN(reset), .Q(LLL4[10]) );
  DFFRHQX1 \LLL5_reg[10]  ( .D(n1000), .CK(clk), .RN(reset), .Q(LLL5[10]) );
  DFFRHQX1 \LLL6_reg[10]  ( .D(n999), .CK(clk), .RN(reset), .Q(LLL6[10]) );
  DFFRHQX1 \LLL2_reg[11]  ( .D(n993), .CK(clk), .RN(reset), .Q(LLL2[11]) );
  DFFRHQX1 \LLL3_reg[11]  ( .D(n992), .CK(clk), .RN(reset), .Q(LLL3[11]) );
  DFFRHQX1 \LLL4_reg[11]  ( .D(n991), .CK(clk), .RN(reset), .Q(LLL4[11]) );
  DFFRHQX1 \LLL5_reg[11]  ( .D(n990), .CK(clk), .RN(reset), .Q(LLL5[11]) );
  DFFRHQX1 \LLL6_reg[11]  ( .D(n989), .CK(clk), .RN(reset), .Q(LLL6[11]) );
  DFFRHQX1 \LLL2_reg[12]  ( .D(n983), .CK(clk), .RN(reset), .Q(LLL2[12]) );
  DFFRHQX1 \LLL3_reg[12]  ( .D(n982), .CK(clk), .RN(reset), .Q(LLL3[12]) );
  DFFRHQX1 \LLL4_reg[12]  ( .D(n981), .CK(clk), .RN(reset), .Q(LLL4[12]) );
  DFFRHQX1 \LLL5_reg[12]  ( .D(n980), .CK(clk), .RN(reset), .Q(LLL5[12]) );
  DFFRHQX1 \LLL6_reg[12]  ( .D(n979), .CK(clk), .RN(reset), .Q(LLL6[12]) );
  DFFRHQX1 \Q2_reg[0]  ( .D(n973), .CK(clk), .RN(reset), .Q(Q2[0]) );
  DFFRHQX1 \Q3_reg[0]  ( .D(n972), .CK(clk), .RN(reset), .Q(Q3[0]) );
  DFFRHQX1 \Q4_reg[0]  ( .D(n971), .CK(clk), .RN(reset), .Q(Q4[0]) );
  DFFRHQX1 \Q5_reg[0]  ( .D(n970), .CK(clk), .RN(reset), .Q(Q5[0]) );
  DFFRHQX1 \Q6_reg[0]  ( .D(n969), .CK(clk), .RN(reset), .Q(Q6[0]) );
  DFFRHQX1 \Q7_reg[0]  ( .D(n968), .CK(clk), .RN(reset), .Q(Q7[0]) );
  DFFRHQX1 \Q2_reg[1]  ( .D(n965), .CK(clk), .RN(reset), .Q(Q2[1]) );
  DFFRHQX1 \Q3_reg[1]  ( .D(n964), .CK(clk), .RN(reset), .Q(Q3[1]) );
  DFFRHQX1 \Q4_reg[1]  ( .D(n963), .CK(clk), .RN(reset), .Q(Q4[1]) );
  DFFRHQX1 \Q5_reg[1]  ( .D(n962), .CK(clk), .RN(reset), .Q(Q5[1]) );
  DFFRHQX1 \Q6_reg[1]  ( .D(n961), .CK(clk), .RN(reset), .Q(Q6[1]) );
  DFFRHQX1 \Q7_reg[1]  ( .D(n960), .CK(clk), .RN(reset), .Q(Q7[1]) );
  DFFRHQX1 \Q2_reg[2]  ( .D(n957), .CK(clk), .RN(reset), .Q(Q2[2]) );
  DFFRHQX1 \Q3_reg[2]  ( .D(n956), .CK(clk), .RN(reset), .Q(Q3[2]) );
  DFFRHQX1 \Q4_reg[2]  ( .D(n955), .CK(clk), .RN(reset), .Q(Q4[2]) );
  DFFRHQX1 \Q5_reg[2]  ( .D(n954), .CK(clk), .RN(reset), .Q(Q5[2]) );
  DFFRHQX1 \Q6_reg[2]  ( .D(n953), .CK(clk), .RN(reset), .Q(Q6[2]) );
  DFFRHQX1 \Q7_reg[2]  ( .D(n952), .CK(clk), .RN(reset), .Q(Q7[2]) );
  DFFRHQX1 \Q2_reg[3]  ( .D(n949), .CK(clk), .RN(reset), .Q(Q2[3]) );
  DFFRHQX1 \Q3_reg[3]  ( .D(n948), .CK(clk), .RN(reset), .Q(Q3[3]) );
  DFFRHQX1 \Q4_reg[3]  ( .D(n947), .CK(clk), .RN(reset), .Q(Q4[3]) );
  DFFRHQX1 \Q5_reg[3]  ( .D(n946), .CK(clk), .RN(reset), .Q(Q5[3]) );
  DFFRHQX1 \Q6_reg[3]  ( .D(n945), .CK(clk), .RN(reset), .Q(Q6[3]) );
  DFFRHQX1 \Q7_reg[3]  ( .D(n944), .CK(clk), .RN(reset), .Q(Q7[3]) );
  DFFRHQX1 \Q2_reg[4]  ( .D(n941), .CK(clk), .RN(reset), .Q(Q2[4]) );
  DFFRHQX1 \Q3_reg[4]  ( .D(n940), .CK(clk), .RN(reset), .Q(Q3[4]) );
  DFFRHQX1 \Q4_reg[4]  ( .D(n939), .CK(clk), .RN(reset), .Q(Q4[4]) );
  DFFRHQX1 \Q5_reg[4]  ( .D(n938), .CK(clk), .RN(reset), .Q(Q5[4]) );
  DFFRHQX1 \Q6_reg[4]  ( .D(n937), .CK(clk), .RN(reset), .Q(Q6[4]) );
  DFFRHQX1 \Q7_reg[4]  ( .D(n936), .CK(clk), .RN(reset), .Q(Q7[4]) );
  DFFRHQX1 \Q2_reg[5]  ( .D(n933), .CK(clk), .RN(reset), .Q(Q2[5]) );
  DFFRHQX1 \Q3_reg[5]  ( .D(n932), .CK(clk), .RN(reset), .Q(Q3[5]) );
  DFFRHQX1 \Q4_reg[5]  ( .D(n931), .CK(clk), .RN(reset), .Q(Q4[5]) );
  DFFRHQX1 \Q5_reg[5]  ( .D(n930), .CK(clk), .RN(reset), .Q(Q5[5]) );
  DFFRHQX1 \Q6_reg[5]  ( .D(n929), .CK(clk), .RN(reset), .Q(Q6[5]) );
  DFFRHQX1 \Q7_reg[5]  ( .D(n928), .CK(clk), .RN(reset), .Q(Q7[5]) );
  DFFRHQX1 \Q2_reg[6]  ( .D(n925), .CK(clk), .RN(reset), .Q(Q2[6]) );
  DFFRHQX1 \Q3_reg[6]  ( .D(n924), .CK(clk), .RN(reset), .Q(Q3[6]) );
  DFFRHQX1 \Q4_reg[6]  ( .D(n923), .CK(clk), .RN(reset), .Q(Q4[6]) );
  DFFRHQX1 \Q5_reg[6]  ( .D(n922), .CK(clk), .RN(reset), .Q(Q5[6]) );
  DFFRHQX1 \Q6_reg[6]  ( .D(n921), .CK(clk), .RN(reset), .Q(Q6[6]) );
  DFFRHQX1 \Q7_reg[6]  ( .D(n920), .CK(clk), .RN(reset), .Q(Q7[6]) );
  DFFRHQX1 \Q2_reg[7]  ( .D(n917), .CK(clk), .RN(reset), .Q(Q2[7]) );
  DFFRHQX1 \Q3_reg[7]  ( .D(n916), .CK(clk), .RN(reset), .Q(Q3[7]) );
  DFFRHQX1 \Q4_reg[7]  ( .D(n915), .CK(clk), .RN(reset), .Q(Q4[7]) );
  DFFRHQX1 \Q5_reg[7]  ( .D(n914), .CK(clk), .RN(reset), .Q(Q5[7]) );
  DFFRHQX1 \Q6_reg[7]  ( .D(n913), .CK(clk), .RN(reset), .Q(Q6[7]) );
  DFFRHQX1 \Q7_reg[7]  ( .D(n912), .CK(clk), .RN(reset), .Q(Q7[7]) );
  DFFRHQX1 \Q2_reg[8]  ( .D(n909), .CK(clk), .RN(reset), .Q(Q2[8]) );
  DFFRHQX1 \Q3_reg[8]  ( .D(n908), .CK(clk), .RN(reset), .Q(Q3[8]) );
  DFFRHQX1 \Q4_reg[8]  ( .D(n907), .CK(clk), .RN(reset), .Q(Q4[8]) );
  DFFRHQX1 \Q5_reg[8]  ( .D(n906), .CK(clk), .RN(reset), .Q(Q5[8]) );
  DFFRHQX1 \Q6_reg[8]  ( .D(n905), .CK(clk), .RN(reset), .Q(Q6[8]) );
  DFFRHQX1 \Q7_reg[8]  ( .D(n904), .CK(clk), .RN(reset), .Q(Q7[8]) );
  DFFRHQX1 \Q2_reg[9]  ( .D(n901), .CK(clk), .RN(reset), .Q(Q2[9]) );
  DFFRHQX1 \Q3_reg[9]  ( .D(n900), .CK(clk), .RN(reset), .Q(Q3[9]) );
  DFFRHQX1 \Q4_reg[9]  ( .D(n899), .CK(clk), .RN(reset), .Q(Q4[9]) );
  DFFRHQX1 \Q5_reg[9]  ( .D(n898), .CK(clk), .RN(reset), .Q(Q5[9]) );
  DFFRHQX1 \Q6_reg[9]  ( .D(n897), .CK(clk), .RN(reset), .Q(Q6[9]) );
  DFFRHQX1 \Q7_reg[9]  ( .D(n896), .CK(clk), .RN(reset), .Q(Q7[9]) );
  DFFRHQX1 \Q2_reg[10]  ( .D(n893), .CK(clk), .RN(reset), .Q(Q2[10]) );
  DFFRHQX1 \Q3_reg[10]  ( .D(n892), .CK(clk), .RN(reset), .Q(Q3[10]) );
  DFFRHQX1 \Q4_reg[10]  ( .D(n891), .CK(clk), .RN(reset), .Q(Q4[10]) );
  DFFRHQX1 \Q5_reg[10]  ( .D(n890), .CK(clk), .RN(reset), .Q(Q5[10]) );
  DFFRHQX1 \Q6_reg[10]  ( .D(n889), .CK(clk), .RN(reset), .Q(Q6[10]) );
  DFFRHQX1 \Q7_reg[10]  ( .D(n888), .CK(clk), .RN(reset), .Q(Q7[10]) );
  DFFRHQX1 \Q2_reg[11]  ( .D(n885), .CK(clk), .RN(reset), .Q(Q2[11]) );
  DFFRHQX1 \Q3_reg[11]  ( .D(n884), .CK(clk), .RN(reset), .Q(Q3[11]) );
  DFFRHQX1 \Q4_reg[11]  ( .D(n883), .CK(clk), .RN(reset), .Q(Q4[11]) );
  DFFRHQX1 \Q5_reg[11]  ( .D(n882), .CK(clk), .RN(reset), .Q(Q5[11]) );
  DFFRHQX1 \Q6_reg[11]  ( .D(n881), .CK(clk), .RN(reset), .Q(Q6[11]) );
  DFFRHQX1 \Q7_reg[11]  ( .D(n880), .CK(clk), .RN(reset), .Q(Q7[11]) );
  DFFRHQX1 \Q2_reg[12]  ( .D(n877), .CK(clk), .RN(reset), .Q(Q2[12]) );
  DFFRHQX1 \Q3_reg[12]  ( .D(n876), .CK(clk), .RN(reset), .Q(Q3[12]) );
  DFFRHQX1 \Q4_reg[12]  ( .D(n875), .CK(clk), .RN(reset), .Q(Q4[12]) );
  DFFRHQX1 \Q5_reg[12]  ( .D(n874), .CK(clk), .RN(reset), .Q(Q5[12]) );
  DFFRHQX1 \Q6_reg[12]  ( .D(n873), .CK(clk), .RN(reset), .Q(Q6[12]) );
  DFFRHQX1 \Q7_reg[12]  ( .D(n872), .CK(clk), .RN(reset), .Q(Q7[12]) );
  DFFRHQX1 \R2_reg[0]  ( .D(n869), .CK(clk), .RN(reset), .Q(R2[0]) );
  DFFRHQX1 \R3_reg[0]  ( .D(n868), .CK(clk), .RN(reset), .Q(R3[0]) );
  DFFRHQX1 \R4_reg[0]  ( .D(n867), .CK(clk), .RN(reset), .Q(R4[0]) );
  DFFRHQX1 \R5_reg[0]  ( .D(n866), .CK(clk), .RN(reset), .Q(R5[0]) );
  DFFRHQX1 \R6_reg[0]  ( .D(n865), .CK(clk), .RN(reset), .Q(R6[0]) );
  DFFRHQX1 \R7_reg[0]  ( .D(n864), .CK(clk), .RN(reset), .Q(R7[0]) );
  DFFRHQX1 \R2_reg[1]  ( .D(n861), .CK(clk), .RN(reset), .Q(R2[1]) );
  DFFRHQX1 \R3_reg[1]  ( .D(n860), .CK(clk), .RN(reset), .Q(R3[1]) );
  DFFRHQX1 \R4_reg[1]  ( .D(n859), .CK(clk), .RN(reset), .Q(R4[1]) );
  DFFRHQX1 \R5_reg[1]  ( .D(n858), .CK(clk), .RN(reset), .Q(R5[1]) );
  DFFRHQX1 \R6_reg[1]  ( .D(n857), .CK(clk), .RN(reset), .Q(R6[1]) );
  DFFRHQX1 \R7_reg[1]  ( .D(n856), .CK(clk), .RN(reset), .Q(R7[1]) );
  DFFRHQX1 \R2_reg[2]  ( .D(n853), .CK(clk), .RN(reset), .Q(R2[2]) );
  DFFRHQX1 \R3_reg[2]  ( .D(n852), .CK(clk), .RN(reset), .Q(R3[2]) );
  DFFRHQX1 \R4_reg[2]  ( .D(n851), .CK(clk), .RN(reset), .Q(R4[2]) );
  DFFRHQX1 \R5_reg[2]  ( .D(n850), .CK(clk), .RN(reset), .Q(R5[2]) );
  DFFRHQX1 \R6_reg[2]  ( .D(n849), .CK(clk), .RN(reset), .Q(R6[2]) );
  DFFRHQX1 \R7_reg[2]  ( .D(n848), .CK(clk), .RN(reset), .Q(R7[2]) );
  DFFRHQX1 \R2_reg[3]  ( .D(n845), .CK(clk), .RN(reset), .Q(R2[3]) );
  DFFRHQX1 \R3_reg[3]  ( .D(n844), .CK(clk), .RN(reset), .Q(R3[3]) );
  DFFRHQX1 \R4_reg[3]  ( .D(n843), .CK(clk), .RN(reset), .Q(R4[3]) );
  DFFRHQX1 \R5_reg[3]  ( .D(n842), .CK(clk), .RN(reset), .Q(R5[3]) );
  DFFRHQX1 \R6_reg[3]  ( .D(n841), .CK(clk), .RN(reset), .Q(R6[3]) );
  DFFRHQX1 \R7_reg[3]  ( .D(n840), .CK(clk), .RN(reset), .Q(R7[3]) );
  DFFRHQX1 \R2_reg[4]  ( .D(n837), .CK(clk), .RN(reset), .Q(R2[4]) );
  DFFRHQX1 \R3_reg[4]  ( .D(n836), .CK(clk), .RN(reset), .Q(R3[4]) );
  DFFRHQX1 \R4_reg[4]  ( .D(n835), .CK(clk), .RN(reset), .Q(R4[4]) );
  DFFRHQX1 \R5_reg[4]  ( .D(n834), .CK(clk), .RN(reset), .Q(R5[4]) );
  DFFRHQX1 \R6_reg[4]  ( .D(n833), .CK(clk), .RN(reset), .Q(R6[4]) );
  DFFRHQX1 \R7_reg[4]  ( .D(n832), .CK(clk), .RN(reset), .Q(R7[4]) );
  DFFRHQX1 \R2_reg[5]  ( .D(n829), .CK(clk), .RN(reset), .Q(R2[5]) );
  DFFRHQX1 \R3_reg[5]  ( .D(n828), .CK(clk), .RN(reset), .Q(R3[5]) );
  DFFRHQX1 \R4_reg[5]  ( .D(n827), .CK(clk), .RN(reset), .Q(R4[5]) );
  DFFRHQX1 \R5_reg[5]  ( .D(n826), .CK(clk), .RN(reset), .Q(R5[5]) );
  DFFRHQX1 \R6_reg[5]  ( .D(n825), .CK(clk), .RN(reset), .Q(R6[5]) );
  DFFRHQX1 \R7_reg[5]  ( .D(n824), .CK(clk), .RN(reset), .Q(R7[5]) );
  DFFRHQX1 \R2_reg[6]  ( .D(n821), .CK(clk), .RN(reset), .Q(R2[6]) );
  DFFRHQX1 \R3_reg[6]  ( .D(n820), .CK(clk), .RN(reset), .Q(R3[6]) );
  DFFRHQX1 \R4_reg[6]  ( .D(n819), .CK(clk), .RN(reset), .Q(R4[6]) );
  DFFRHQX1 \R5_reg[6]  ( .D(n818), .CK(clk), .RN(reset), .Q(R5[6]) );
  DFFRHQX1 \R6_reg[6]  ( .D(n817), .CK(clk), .RN(reset), .Q(R6[6]) );
  DFFRHQX1 \R7_reg[6]  ( .D(n816), .CK(clk), .RN(reset), .Q(R7[6]) );
  DFFRHQX1 \R2_reg[7]  ( .D(n813), .CK(clk), .RN(reset), .Q(R2[7]) );
  DFFRHQX1 \R3_reg[7]  ( .D(n812), .CK(clk), .RN(reset), .Q(R3[7]) );
  DFFRHQX1 \R4_reg[7]  ( .D(n811), .CK(clk), .RN(reset), .Q(R4[7]) );
  DFFRHQX1 \R5_reg[7]  ( .D(n810), .CK(clk), .RN(reset), .Q(R5[7]) );
  DFFRHQX1 \R6_reg[7]  ( .D(n809), .CK(clk), .RN(reset), .Q(R6[7]) );
  DFFRHQX1 \R7_reg[7]  ( .D(n808), .CK(clk), .RN(reset), .Q(R7[7]) );
  DFFRHQX1 \R2_reg[8]  ( .D(n805), .CK(clk), .RN(reset), .Q(R2[8]) );
  DFFRHQX1 \R3_reg[8]  ( .D(n804), .CK(clk), .RN(reset), .Q(R3[8]) );
  DFFRHQX1 \R4_reg[8]  ( .D(n803), .CK(clk), .RN(reset), .Q(R4[8]) );
  DFFRHQX1 \R5_reg[8]  ( .D(n802), .CK(clk), .RN(reset), .Q(R5[8]) );
  DFFRHQX1 \R6_reg[8]  ( .D(n801), .CK(clk), .RN(reset), .Q(R6[8]) );
  DFFRHQX1 \R7_reg[8]  ( .D(n800), .CK(clk), .RN(reset), .Q(R7[8]) );
  DFFRHQX1 \R2_reg[9]  ( .D(n797), .CK(clk), .RN(reset), .Q(R2[9]) );
  DFFRHQX1 \R3_reg[9]  ( .D(n796), .CK(clk), .RN(reset), .Q(R3[9]) );
  DFFRHQX1 \R4_reg[9]  ( .D(n795), .CK(clk), .RN(reset), .Q(R4[9]) );
  DFFRHQX1 \R5_reg[9]  ( .D(n794), .CK(clk), .RN(reset), .Q(R5[9]) );
  DFFRHQX1 \R6_reg[9]  ( .D(n793), .CK(clk), .RN(reset), .Q(R6[9]) );
  DFFRHQX1 \R7_reg[9]  ( .D(n792), .CK(clk), .RN(reset), .Q(R7[9]) );
  DFFRHQX1 \R2_reg[10]  ( .D(n789), .CK(clk), .RN(reset), .Q(R2[10]) );
  DFFRHQX1 \R3_reg[10]  ( .D(n788), .CK(clk), .RN(reset), .Q(R3[10]) );
  DFFRHQX1 \R4_reg[10]  ( .D(n787), .CK(clk), .RN(reset), .Q(R4[10]) );
  DFFRHQX1 \R5_reg[10]  ( .D(n786), .CK(clk), .RN(reset), .Q(R5[10]) );
  DFFRHQX1 \R6_reg[10]  ( .D(n785), .CK(clk), .RN(reset), .Q(R6[10]) );
  DFFRHQX1 \R7_reg[10]  ( .D(n784), .CK(clk), .RN(reset), .Q(R7[10]) );
  DFFRHQX1 \R2_reg[11]  ( .D(n781), .CK(clk), .RN(reset), .Q(R2[11]) );
  DFFRHQX1 \R3_reg[11]  ( .D(n780), .CK(clk), .RN(reset), .Q(R3[11]) );
  DFFRHQX1 \R4_reg[11]  ( .D(n779), .CK(clk), .RN(reset), .Q(R4[11]) );
  DFFRHQX1 \R5_reg[11]  ( .D(n778), .CK(clk), .RN(reset), .Q(R5[11]) );
  DFFRHQX1 \R6_reg[11]  ( .D(n777), .CK(clk), .RN(reset), .Q(R6[11]) );
  DFFRHQX1 \R7_reg[11]  ( .D(n776), .CK(clk), .RN(reset), .Q(R7[11]) );
  DFFRHQX1 \R2_reg[12]  ( .D(n773), .CK(clk), .RN(reset), .Q(R2[12]) );
  DFFRHQX1 \R3_reg[12]  ( .D(n772), .CK(clk), .RN(reset), .Q(R3[12]) );
  DFFRHQX1 \R4_reg[12]  ( .D(n771), .CK(clk), .RN(reset), .Q(R4[12]) );
  DFFRHQX1 \R5_reg[12]  ( .D(n770), .CK(clk), .RN(reset), .Q(R5[12]) );
  DFFRHQX1 \R6_reg[12]  ( .D(n769), .CK(clk), .RN(reset), .Q(R6[12]) );
  DFFRHQX1 \R7_reg[12]  ( .D(n768), .CK(clk), .RN(reset), .Q(R7[12]) );
  DFFRHQX1 ST1_reg ( .D(n755), .CK(clk), .RN(reset), .Q(ST1) );
  DFFRHQX1 \DQ1_reg[0]  ( .D(n753), .CK(clk), .RN(reset), .Q(DQ1[0]) );
  DFFRHQX1 \DQ2_reg[0]  ( .D(n752), .CK(clk), .RN(reset), .Q(DQ2[0]) );
  DFFRHQX1 \DQ3_reg[0]  ( .D(n751), .CK(clk), .RN(reset), .Q(DQ3[0]) );
  DFFRHQX1 \DQ4_reg[0]  ( .D(n750), .CK(clk), .RN(reset), .Q(DQ4[0]) );
  DFFRHQX1 \DQ5_reg[0]  ( .D(n749), .CK(clk), .RN(reset), .Q(DQ5[0]) );
  DFFRHQX1 \DQ6_reg[0]  ( .D(n748), .CK(clk), .RN(reset), .Q(DQ6[0]) );
  DFFRHQX1 \DQ1_reg[1]  ( .D(n745), .CK(clk), .RN(reset), .Q(DQ1[1]) );
  DFFRHQX1 \DQ2_reg[1]  ( .D(n744), .CK(clk), .RN(reset), .Q(DQ2[1]) );
  DFFRHQX1 \DQ3_reg[1]  ( .D(n743), .CK(clk), .RN(reset), .Q(DQ3[1]) );
  DFFRHQX1 \DQ4_reg[1]  ( .D(n742), .CK(clk), .RN(reset), .Q(DQ4[1]) );
  DFFRHQX1 \DQ5_reg[1]  ( .D(n741), .CK(clk), .RN(reset), .Q(DQ5[1]) );
  DFFRHQX1 \DQ6_reg[1]  ( .D(n740), .CK(clk), .RN(reset), .Q(DQ6[1]) );
  DFFRHQX1 \DQ1_reg[2]  ( .D(n737), .CK(clk), .RN(reset), .Q(DQ1[2]) );
  DFFRHQX1 \DQ2_reg[2]  ( .D(n736), .CK(clk), .RN(reset), .Q(DQ2[2]) );
  DFFRHQX1 \DQ3_reg[2]  ( .D(n735), .CK(clk), .RN(reset), .Q(DQ3[2]) );
  DFFRHQX1 \DQ4_reg[2]  ( .D(n734), .CK(clk), .RN(reset), .Q(DQ4[2]) );
  DFFRHQX1 \DQ5_reg[2]  ( .D(n733), .CK(clk), .RN(reset), .Q(DQ5[2]) );
  DFFRHQX1 \DQ6_reg[2]  ( .D(n732), .CK(clk), .RN(reset), .Q(DQ6[2]) );
  DFFRHQX1 \DQ1_reg[3]  ( .D(n729), .CK(clk), .RN(reset), .Q(DQ1[3]) );
  DFFRHQX1 \DQ2_reg[3]  ( .D(n728), .CK(clk), .RN(reset), .Q(DQ2[3]) );
  DFFRHQX1 \DQ3_reg[3]  ( .D(n727), .CK(clk), .RN(reset), .Q(DQ3[3]) );
  DFFRHQX1 \DQ4_reg[3]  ( .D(n726), .CK(clk), .RN(reset), .Q(DQ4[3]) );
  DFFRHQX1 \DQ5_reg[3]  ( .D(n725), .CK(clk), .RN(reset), .Q(DQ5[3]) );
  DFFRHQX1 \DQ6_reg[3]  ( .D(n724), .CK(clk), .RN(reset), .Q(DQ6[3]) );
  DFFRHQX1 \DQ1_reg[4]  ( .D(n721), .CK(clk), .RN(reset), .Q(DQ1[4]) );
  DFFRHQX1 \DQ2_reg[4]  ( .D(n720), .CK(clk), .RN(reset), .Q(DQ2[4]) );
  DFFRHQX1 \DQ3_reg[4]  ( .D(n719), .CK(clk), .RN(reset), .Q(DQ3[4]) );
  DFFRHQX1 \DQ4_reg[4]  ( .D(n718), .CK(clk), .RN(reset), .Q(DQ4[4]) );
  DFFRHQX1 \DQ5_reg[4]  ( .D(n717), .CK(clk), .RN(reset), .Q(DQ5[4]) );
  DFFRHQX1 \DQ6_reg[4]  ( .D(n716), .CK(clk), .RN(reset), .Q(DQ6[4]) );
  DFFRHQX1 \DR1_reg[0]  ( .D(n713), .CK(clk), .RN(reset), .Q(DR1[0]) );
  DFFRHQX1 \DR2_reg[0]  ( .D(n712), .CK(clk), .RN(reset), .Q(DR2[0]) );
  DFFRHQX1 \DR3_reg[0]  ( .D(n711), .CK(clk), .RN(reset), .Q(DR3[0]) );
  DFFRHQX1 \DR4_reg[0]  ( .D(n710), .CK(clk), .RN(reset), .Q(DR4[0]) );
  DFFRHQX1 \DR5_reg[0]  ( .D(n709), .CK(clk), .RN(reset), .Q(DR5[0]) );
  DFFRHQX1 \DR6_reg[0]  ( .D(n708), .CK(clk), .RN(reset), .Q(DR6[0]) );
  DFFRHQX1 \DR1_reg[1]  ( .D(n705), .CK(clk), .RN(reset), .Q(DR1[1]) );
  DFFRHQX1 \DR2_reg[1]  ( .D(n704), .CK(clk), .RN(reset), .Q(DR2[1]) );
  DFFRHQX1 \DR3_reg[1]  ( .D(n703), .CK(clk), .RN(reset), .Q(DR3[1]) );
  DFFRHQX1 \DR4_reg[1]  ( .D(n702), .CK(clk), .RN(reset), .Q(DR4[1]) );
  DFFRHQX1 \DR5_reg[1]  ( .D(n701), .CK(clk), .RN(reset), .Q(DR5[1]) );
  DFFRHQX1 \DR6_reg[1]  ( .D(n700), .CK(clk), .RN(reset), .Q(DR6[1]) );
  DFFRHQX1 \DR1_reg[2]  ( .D(n697), .CK(clk), .RN(reset), .Q(DR1[2]) );
  DFFRHQX1 \DR2_reg[2]  ( .D(n696), .CK(clk), .RN(reset), .Q(DR2[2]) );
  DFFRHQX1 \DR3_reg[2]  ( .D(n695), .CK(clk), .RN(reset), .Q(DR3[2]) );
  DFFRHQX1 \DR4_reg[2]  ( .D(n694), .CK(clk), .RN(reset), .Q(DR4[2]) );
  DFFRHQX1 \DR5_reg[2]  ( .D(n693), .CK(clk), .RN(reset), .Q(DR5[2]) );
  DFFRHQX1 \DR6_reg[2]  ( .D(n692), .CK(clk), .RN(reset), .Q(DR6[2]) );
  DFFRHQX1 \DR1_reg[3]  ( .D(n689), .CK(clk), .RN(reset), .Q(DR1[3]) );
  DFFRHQX1 \DR2_reg[3]  ( .D(n688), .CK(clk), .RN(reset), .Q(DR2[3]) );
  DFFRHQX1 \DR3_reg[3]  ( .D(n687), .CK(clk), .RN(reset), .Q(DR3[3]) );
  DFFRHQX1 \DR4_reg[3]  ( .D(n686), .CK(clk), .RN(reset), .Q(DR4[3]) );
  DFFRHQX1 \DR5_reg[3]  ( .D(n685), .CK(clk), .RN(reset), .Q(DR5[3]) );
  DFFRHQX1 \DR6_reg[3]  ( .D(n684), .CK(clk), .RN(reset), .Q(DR6[3]) );
  DFFRHQX1 \DR1_reg[4]  ( .D(n681), .CK(clk), .RN(reset), .Q(DR1[4]) );
  DFFRHQX1 \DR2_reg[4]  ( .D(n680), .CK(clk), .RN(reset), .Q(DR2[4]) );
  DFFRHQX1 \DR3_reg[4]  ( .D(n679), .CK(clk), .RN(reset), .Q(DR3[4]) );
  DFFRHQX1 \DR4_reg[4]  ( .D(n678), .CK(clk), .RN(reset), .Q(DR4[4]) );
  DFFRHQX1 \DR5_reg[4]  ( .D(n677), .CK(clk), .RN(reset), .Q(DR5[4]) );
  DFFRHQX1 \DR6_reg[4]  ( .D(n676), .CK(clk), .RN(reset), .Q(DR6[4]) );
  DFFRHQX1 \dR_reg_reg[4]  ( .D(n1313), .CK(clk), .RN(reset), .Q(dR_reg[4]) );
  DFFRHQX1 \dQ_reg_reg[4]  ( .D(n1308), .CK(clk), .RN(reset), .Q(dQ_reg[4]) );
  DFFRHQX1 \Rin_reg_reg[9]  ( .D(n1298), .CK(clk), .RN(reset), .Q(Rin_reg[9])
         );
  DFFRHQX1 \Qin_reg_reg[9]  ( .D(n1285), .CK(clk), .RN(reset), .Q(Qin_reg[9])
         );
  DFFRHQX1 \Uin_reg_reg[9]  ( .D(n1259), .CK(clk), .RN(reset), .Q(Uin_reg[9])
         );
  DFFRHQX1 \count_reg[9]  ( .D(n1240), .CK(clk), .RN(reset), .Q(count[9]) );
  DFFRHQX1 ST2_reg ( .D(n754), .CK(clk), .RN(reset), .Q(ST2) );
  DFFRHQX1 \count_reg[8]  ( .D(n1241), .CK(clk), .RN(reset), .Q(count[8]) );
  DFFRHQX1 \count_reg[7]  ( .D(n1242), .CK(clk), .RN(reset), .Q(count[7]) );
  DFFSX1 \stop1_reg[2]  ( .D(n1236), .CK(clk), .SN(reset), .Q(stop1[2]), .QN(
        n645) );
  DFFSX1 \stop2_reg[2]  ( .D(n1233), .CK(clk), .SN(reset), .Q(stop2[2]), .QN(
        n648) );
  DFFSX1 \s_reg_reg[2]  ( .D(n756), .CK(clk), .SN(reset), .Q(s_reg[2]), .QN(
        n654) );
  DFFRHQX1 \DQ8_reg[3]  ( .D(n722), .CK(clk), .RN(reset), .Q(DQ8[3]) );
  DFFRHQX1 \dQ_reg_reg[3]  ( .D(n1307), .CK(clk), .RN(reset), .Q(dQ_reg[3]) );
  DFFRHQX1 \count_reg[0]  ( .D(n1249), .CK(clk), .RN(reset), .Q(count[0]) );
  DFFRHQX1 \count_reg[2]  ( .D(n1247), .CK(clk), .RN(reset), .Q(count[2]) );
  DFFRHQX1 \count_reg[4]  ( .D(n1245), .CK(clk), .RN(reset), .Q(count[4]) );
  DFFRHQX1 \count_reg[5]  ( .D(n1244), .CK(clk), .RN(reset), .Q(count[5]) );
  DFFRHQX1 \count_reg[1]  ( .D(n1248), .CK(clk), .RN(reset), .Q(count[1]) );
  DFFRHQX1 \count_reg[6]  ( .D(n1243), .CK(clk), .RN(reset), .Q(count[6]) );
  DFFRHQX1 \count_reg[3]  ( .D(n1246), .CK(clk), .RN(reset), .Q(count[3]) );
  DFFSX1 St_reg_reg ( .D(n1303), .CK(clk), .SN(reset), .Q(St_reg), .QN(n673)
         );
  DFFSX1 feedback_sel_reg ( .D(n1239), .CK(clk), .SN(reset), .Q(feedback_sel), 
        .QN(n671) );
  DFFSX1 \stop3_reg[2]  ( .D(n1230), .CK(clk), .SN(reset), .Q(stop3[2]), .QN(
        n651) );
  DFFRHQXL \LLL1_reg[9]  ( .D(n1419), .CK(clk), .RN(reset), .Q(LLL1[9]) );
  DFFRHQXL \LLL1_reg[10]  ( .D(n1421), .CK(clk), .RN(reset), .Q(LLL1[10]) );
  DFFRHQXL \L1_reg[9]  ( .D(n1420), .CK(clk), .RN(reset), .Q(L1[9]) );
  DFFRHQXL \L1_reg[10]  ( .D(n1422), .CK(clk), .RN(reset), .Q(L1[10]) );
  DFFRHQXL \R1_reg[4]  ( .D(n1426), .CK(clk), .RN(reset), .Q(R1[4]) );
  DFFRHQXL \R1_reg[8]  ( .D(n1429), .CK(clk), .RN(reset), .Q(R1[8]) );
  DFFRHQXL \R1_reg[9]  ( .D(n1430), .CK(clk), .RN(reset), .Q(R1[9]) );
  DFFRHQXL \R1_reg[10]  ( .D(n1431), .CK(clk), .RN(reset), .Q(R1[10]) );
  DFFRHQXL \R1_reg[11]  ( .D(n1432), .CK(clk), .RN(reset), .Q(R1[11]) );
  MX2X1 U3_inst ( .A(R1[11]), .B(Rout[11]), .S0(N99), .Y(n1432) );
  MX2X1 U4_inst ( .A(R1[10]), .B(Rout[10]), .S0(n1398), .Y(n1431) );
  MX2X1 U5_inst ( .A(R1[9]), .B(Rout[9]), .S0(n1396), .Y(n1430) );
  MX2X1 U6_inst ( .A(R1[8]), .B(Rout[8]), .S0(n1398), .Y(n1429) );
  MX2X1 U7_inst ( .A(R1[4]), .B(Rout[4]), .S0(n1393), .Y(n1426) );
  INVX1 U8_inst ( .A(R1[12]), .Y(n1) );
  MX2X1 U9 ( .A(R1[7]), .B(Rout[7]), .S0(n1392), .Y(n1428) );
  MX2X1 U10 ( .A(R1[3]), .B(Rout[3]), .S0(n643), .Y(n1425) );
  MX2X1 U11 ( .A(R1[5]), .B(Rout[5]), .S0(n1399), .Y(n1427) );
  MX2X1 U12 ( .A(L1[3]), .B(Lout_temp[3]), .S0(n1394), .Y(n1410) );
  MX2X1 U13 ( .A(Lout_temp[3]), .B(LLL1[3]), .S0(n1383), .Y(n1409) );
  AOI2BB2X1 U14 ( .B0(Rout[12]), .B1(n1046), .A0N(n1393), .A1N(n1), .Y(n106)
         );
  AOI22X1 U15 ( .A0(n650), .A1(Lout_temp[0]), .B0(n1356), .B1(LLL1[0]), .Y(
        n436) );
  INVXL U16 ( .A(n106), .Y(n774) );
  INVXL U17 ( .A(n308), .Y(n976) );
  INVXL U18 ( .A(n316), .Y(n984) );
  INVXL U19 ( .A(n186), .Y(n854) );
  INVXL U20 ( .A(n154), .Y(n822) );
  INVXL U21 ( .A(n194), .Y(n862) );
  INVXL U22 ( .A(n368), .Y(n1036) );
  INVXL U23 ( .A(n376), .Y(n1044) );
  INVXL U24 ( .A(n428), .Y(n1096) );
  INVXL U25 ( .A(n436), .Y(n1104) );
  INVXL U26 ( .A(n418), .Y(n1086) );
  INVXL U27 ( .A(n426), .Y(n1094) );
  INVXL U28 ( .A(n408), .Y(n1076) );
  INVXL U29 ( .A(n416), .Y(n1084) );
  INVX1 U30 ( .A(n1381), .Y(n814) );
  INVX1 U31 ( .A(n1381), .Y(n830) );
  INVX1 U32 ( .A(n1381), .Y(n838) );
  INVX1 U33 ( .A(n1380), .Y(n846) );
  INVX1 U34 ( .A(n1380), .Y(n986) );
  INVX1 U35 ( .A(n1380), .Y(n994) );
  INVX1 U36 ( .A(n1379), .Y(n996) );
  INVX1 U37 ( .A(n1377), .Y(n1026) );
  INVX1 U38 ( .A(n1377), .Y(n1024) );
  INVX1 U39 ( .A(n1378), .Y(n1016) );
  INVX1 U40 ( .A(n1378), .Y(n1006) );
  INVX1 U41 ( .A(n1378), .Y(n1014) );
  INVX1 U42 ( .A(n1386), .Y(n661) );
  INVX1 U43 ( .A(n1386), .Y(n660) );
  INVX1 U44 ( .A(n1386), .Y(n659) );
  INVX1 U45 ( .A(n1387), .Y(n658) );
  INVX1 U46 ( .A(n1387), .Y(n657) );
  INVX1 U47 ( .A(n1387), .Y(n656) );
  INVX1 U48 ( .A(n1382), .Y(n806) );
  INVX1 U49 ( .A(n1382), .Y(n798) );
  INVX1 U50 ( .A(n1382), .Y(n790) );
  INVX1 U51 ( .A(n1383), .Y(n782) );
  INVX1 U52 ( .A(n1379), .Y(n1004) );
  INVX1 U53 ( .A(n1383), .Y(n670) );
  INVX1 U54 ( .A(n1383), .Y(n669) );
  INVX1 U55 ( .A(n1384), .Y(n667) );
  INVX1 U56 ( .A(n1384), .Y(n666) );
  INVX1 U57 ( .A(n1385), .Y(n665) );
  INVX1 U58 ( .A(n1385), .Y(n664) );
  INVX1 U59 ( .A(n1385), .Y(n662) );
  INVX1 U60 ( .A(n1384), .Y(n668) );
  INVX1 U61 ( .A(n1377), .Y(n1034) );
  INVX1 U62 ( .A(n1376), .Y(n1054) );
  INVX1 U63 ( .A(n1376), .Y(n1056) );
  INVX1 U64 ( .A(n1375), .Y(n1064) );
  INVX1 U65 ( .A(n1375), .Y(n1066) );
  INVX1 U66 ( .A(n1375), .Y(n1074) );
  INVX1 U67 ( .A(n1374), .Y(n1314) );
  INVX1 U68 ( .A(n1374), .Y(n1315) );
  INVX1 U69 ( .A(n1376), .Y(n1046) );
  INVX1 U70 ( .A(n1374), .Y(n1316) );
  INVX1 U71 ( .A(n1373), .Y(n1318) );
  INVX1 U72 ( .A(n1373), .Y(n1319) );
  INVX1 U73 ( .A(n1373), .Y(n1317) );
  INVX1 U74 ( .A(n1372), .Y(n1321) );
  INVX1 U75 ( .A(n1372), .Y(n1322) );
  INVX1 U76 ( .A(n1371), .Y(n1323) );
  INVX1 U77 ( .A(n1371), .Y(n1324) );
  INVX1 U78 ( .A(n1371), .Y(n1325) );
  INVX1 U79 ( .A(n1372), .Y(n1320) );
  INVX1 U80 ( .A(n1370), .Y(n1328) );
  INVX1 U81 ( .A(n1370), .Y(n1326) );
  INVX1 U82 ( .A(n1370), .Y(n1327) );
  INVX1 U83 ( .A(n1379), .Y(n1329) );
  INVX1 U84 ( .A(n643), .Y(n1335) );
  INVX1 U85 ( .A(n1399), .Y(n1333) );
  INVX1 U86 ( .A(n1397), .Y(n1334) );
  INVX1 U87 ( .A(n643), .Y(n1331) );
  INVX1 U88 ( .A(n1396), .Y(n1330) );
  INVX1 U89 ( .A(n1395), .Y(n1332) );
  INVX1 U90 ( .A(n643), .Y(n1338) );
  INVX1 U91 ( .A(n1398), .Y(n1336) );
  INVX1 U92 ( .A(n1395), .Y(n1337) );
  INVX1 U93 ( .A(n1395), .Y(n1339) );
  INVX1 U94 ( .A(n1397), .Y(n1340) );
  INVX1 U95 ( .A(n1394), .Y(n1341) );
  INVX1 U96 ( .A(n1391), .Y(n1348) );
  INVX1 U97 ( .A(n643), .Y(n1346) );
  INVX1 U98 ( .A(n1399), .Y(n1366) );
  INVX1 U99 ( .A(n643), .Y(n1343) );
  INVX1 U100 ( .A(n1399), .Y(n1342) );
  INVX1 U101 ( .A(N99), .Y(n1345) );
  INVX1 U102 ( .A(n1399), .Y(n1353) );
  INVX1 U103 ( .A(n1399), .Y(n1344) );
  INVX1 U104 ( .A(n1396), .Y(n1347) );
  INVX1 U105 ( .A(n643), .Y(n1361) );
  INVX1 U106 ( .A(n1396), .Y(n1351) );
  INVX1 U107 ( .A(n1399), .Y(n1350) );
  INVX1 U108 ( .A(n1398), .Y(n1349) );
  INVX1 U109 ( .A(n644), .Y(n1352) );
  INVX1 U110 ( .A(n1394), .Y(n1354) );
  INVX1 U111 ( .A(n1391), .Y(n1359) );
  INVX1 U112 ( .A(n1398), .Y(n1368) );
  INVX1 U113 ( .A(n1392), .Y(n1356) );
  INVX1 U114 ( .A(n1393), .Y(n1355) );
  INVX1 U115 ( .A(n1397), .Y(n1357) );
  INVX1 U116 ( .A(n1398), .Y(n1362) );
  INVX1 U117 ( .A(n643), .Y(n1358) );
  INVX1 U118 ( .A(n643), .Y(n1360) );
  INVX1 U119 ( .A(n1399), .Y(n1364) );
  INVX1 U120 ( .A(n1398), .Y(n1363) );
  INVX1 U121 ( .A(n1398), .Y(n1367) );
  INVX1 U122 ( .A(n1399), .Y(n1365) );
  INVX1 U123 ( .A(n1398), .Y(n1369) );
  INVX1 U124 ( .A(n1390), .Y(n644) );
  INVX1 U125 ( .A(n1390), .Y(n643) );
  INVX1 U126 ( .A(n1390), .Y(n646) );
  INVX1 U127 ( .A(n1389), .Y(n647) );
  INVX1 U128 ( .A(n1389), .Y(n649) );
  INVX1 U129 ( .A(n1388), .Y(n653) );
  INVX1 U130 ( .A(n1388), .Y(n652) );
  INVX1 U131 ( .A(n1389), .Y(n650) );
  INVX1 U132 ( .A(n1388), .Y(n655) );
  INVX1 U133 ( .A(n1396), .Y(n1373) );
  INVX1 U134 ( .A(n1394), .Y(n1381) );
  INVX1 U135 ( .A(n1394), .Y(n1380) );
  INVX1 U136 ( .A(n1395), .Y(n1377) );
  INVX1 U137 ( .A(n1395), .Y(n1378) );
  INVX1 U138 ( .A(n1392), .Y(n1386) );
  INVX1 U139 ( .A(n1397), .Y(n1371) );
  INVX1 U140 ( .A(n1397), .Y(n1372) );
  INVX1 U141 ( .A(n1397), .Y(n1370) );
  INVX1 U142 ( .A(n1392), .Y(n1387) );
  INVX1 U143 ( .A(n1393), .Y(n1382) );
  INVX1 U144 ( .A(n1394), .Y(n1379) );
  INVX1 U145 ( .A(n1393), .Y(n1383) );
  INVX1 U146 ( .A(n1392), .Y(n1385) );
  INVX1 U147 ( .A(n1393), .Y(n1384) );
  INVX1 U148 ( .A(n1403), .Y(n1399) );
  INVX1 U149 ( .A(n1403), .Y(n1398) );
  INVX1 U150 ( .A(n1396), .Y(n1375) );
  INVX1 U151 ( .A(n1396), .Y(n1374) );
  INVX1 U152 ( .A(n1395), .Y(n1376) );
  INVX1 U153 ( .A(n1391), .Y(n1390) );
  INVX1 U154 ( .A(n1396), .Y(n1401) );
  INVX1 U155 ( .A(n1404), .Y(n1397) );
  INVX1 U156 ( .A(n1405), .Y(n1394) );
  INVX1 U157 ( .A(n1405), .Y(n1392) );
  INVX1 U158 ( .A(n1405), .Y(n1393) );
  INVX1 U159 ( .A(n1392), .Y(n1400) );
  INVX1 U160 ( .A(n1395), .Y(n1402) );
  INVX1 U161 ( .A(n1395), .Y(n1403) );
  INVX1 U162 ( .A(n1404), .Y(n1396) );
  INVX1 U163 ( .A(n1404), .Y(n1395) );
  INVX1 U164 ( .A(n1391), .Y(n1388) );
  INVX1 U165 ( .A(n1391), .Y(n1389) );
  INVX1 U166 ( .A(n1406), .Y(n1391) );
  INVX1 U167 ( .A(n1407), .Y(n1406) );
  INVX1 U168 ( .A(n1407), .Y(n1405) );
  INVX1 U169 ( .A(n1407), .Y(n1404) );
  INVX1 U170 ( .A(n1408), .Y(n1407) );
  INVX1 U171 ( .A(n671), .Y(n406) );
  INVX1 U172 ( .A(n671), .Y(n398) );
  INVX1 U173 ( .A(n562), .Y(n1232) );
  AOI22X1 U174 ( .A0(n1334), .A1(stop3[0]), .B0(Lstop3), .B1(n1056), .Y(n562)
         );
  INVX1 U175 ( .A(n564), .Y(n1235) );
  AOI22X1 U176 ( .A0(n1340), .A1(stop2[0]), .B0(Lstop2), .B1(n1056), .Y(n564)
         );
  INVX1 U177 ( .A(n566), .Y(n1238) );
  AOI22X1 U178 ( .A0(n1359), .A1(stop1[0]), .B0(Lstop1), .B1(n1056), .Y(n566)
         );
  MX2X1 U179 ( .A(LLL1[4]), .B(Lout_temp[4]), .S0(N99), .Y(n1411) );
  MX2X1 U180 ( .A(L1[4]), .B(Lout_temp[4]), .S0(n1393), .Y(n1412) );
  AOI22X1 U181 ( .A0(n655), .A1(Lout_temp[12]), .B0(n1362), .B1(L1[12]), .Y(
        n308) );
  MX2X1 U182 ( .A(L1[8]), .B(Lout_temp[8]), .S0(n1398), .Y(n1418) );
  MX2X1 U183 ( .A(LLL1[8]), .B(Lout_temp[8]), .S0(n1392), .Y(n1417) );
  MX2X1 U184 ( .A(L1[7]), .B(Lout_temp[7]), .S0(n1397), .Y(n1416) );
  MX2X1 U185 ( .A(LLL1[7]), .B(Lout_temp[7]), .S0(n1396), .Y(n1415) );
  MX2X1 U186 ( .A(L1[5]), .B(Lout_temp[5]), .S0(n1394), .Y(n1414) );
  MX2X1 U187 ( .A(LLL1[5]), .B(Lout_temp[5]), .S0(n1397), .Y(n1413) );
  MX2X1 U188 ( .A(L1[11]), .B(Lout_temp[11]), .S0(N99), .Y(n1424) );
  MX2X1 U189 ( .A(LLL1[11]), .B(Lout_temp[11]), .S0(n1394), .Y(n1423) );
  MX2X1 U190 ( .A(L1[10]), .B(Lout_temp[10]), .S0(n1393), .Y(n1422) );
  MX2X1 U191 ( .A(LLL1[10]), .B(Lout_temp[10]), .S0(n1395), .Y(n1421) );
  MX2X1 U192 ( .A(L1[9]), .B(Lout_temp[9]), .S0(n1392), .Y(n1420) );
  MX2X1 U193 ( .A(LLL1[9]), .B(Lout_temp[9]), .S0(n1393), .Y(n1419) );
  AOI22X1 U194 ( .A0(n655), .A1(Lout_temp[12]), .B0(n1363), .B1(LLL1[12]), .Y(
        n316) );
  AOI22X1 U195 ( .A0(n653), .A1(Lout_temp[6]), .B0(n1362), .B1(L1[6]), .Y(n368) );
  AOI22X1 U196 ( .A0(n653), .A1(Lout_temp[6]), .B0(n1390), .B1(LLL1[6]), .Y(
        n376) );
  AOI22X1 U197 ( .A0(n652), .A1(Lout_temp[2]), .B0(n1334), .B1(L1[2]), .Y(n408) );
  AOI22X1 U198 ( .A0(n652), .A1(Lout_temp[2]), .B0(n1339), .B1(LLL1[2]), .Y(
        n416) );
  AOI22X1 U199 ( .A0(n650), .A1(Lout_temp[1]), .B0(n1372), .B1(L1[1]), .Y(n418) );
  AOI22X1 U200 ( .A0(n650), .A1(Lout_temp[1]), .B0(n1390), .B1(LLL1[1]), .Y(
        n426) );
  AOI22X1 U201 ( .A0(n650), .A1(Lout_temp[0]), .B0(n1360), .B1(L1[0]), .Y(n428) );
  INVX1 U202 ( .A(n88), .Y(n755) );
  AOI22X1 U203 ( .A0(n814), .A1(stop_o), .B0(n1340), .B1(ST1), .Y(n88) );
  INVX1 U204 ( .A(n525), .Y(n1193) );
  AOI22X1 U205 ( .A0(n666), .A1(Uout[3]), .B0(n1355), .B1(U1[3]), .Y(n525) );
  INVX1 U206 ( .A(n534), .Y(n1202) );
  AOI22X1 U207 ( .A0(n666), .A1(Uout[2]), .B0(n1388), .B1(U1[2]), .Y(n534) );
  AOI22X1 U208 ( .A0(n1357), .A1(R1[6]), .B0(Rout[6]), .B1(n1074), .Y(n154) );
  AOI22X1 U209 ( .A0(n1336), .A1(R1[2]), .B0(Rout[2]), .B1(n1054), .Y(n186) );
  AOI22X1 U210 ( .A0(n1337), .A1(R1[1]), .B0(Rout[1]), .B1(n1046), .Y(n194) );
  INVX1 U211 ( .A(n202), .Y(n870) );
  AOI22X1 U212 ( .A0(n1360), .A1(R1[0]), .B0(Rout[0]), .B1(n1054), .Y(n202) );
  INVX1 U213 ( .A(n526), .Y(n1194) );
  AOI22X1 U214 ( .A0(n666), .A1(Uout[3]), .B0(Uout_temp[3]), .B1(n1341), .Y(
        n526) );
  INVX1 U215 ( .A(n535), .Y(n1203) );
  AOI22X1 U216 ( .A0(n665), .A1(Uout[2]), .B0(Uout_temp[2]), .B1(n1400), .Y(
        n535) );
  INVX1 U217 ( .A(n98), .Y(n766) );
  AOI22X1 U218 ( .A0(n830), .A1(stop_o), .B0(n1384), .B1(STOP1), .Y(n98) );
  NOR4X1 U219 ( .A(out_sel[9]), .B(out_sel[8]), .C(out_sel[7]), .D(out_sel[6]), 
        .Y(n5) );
  NOR3X1 U220 ( .A(out_sel[3]), .B(out_sel[5]), .C(out_sel[4]), .Y(n4) );
  INVX1 U221 ( .A(n90), .Y(n758) );
  AOI22X1 U222 ( .A0(n814), .A1(STOP8), .B0(n1382), .B1(s_reg[0]), .Y(n90) );
  INVX1 U223 ( .A(n91), .Y(n759) );
  AOI22X1 U224 ( .A0(n814), .A1(STOP7), .B0(n1385), .B1(STOP8), .Y(n91) );
  INVX1 U225 ( .A(n92), .Y(n760) );
  AOI22X1 U226 ( .A0(n814), .A1(STOP6), .B0(n1364), .B1(STOP7), .Y(n92) );
  INVX1 U227 ( .A(n93), .Y(n761) );
  AOI22X1 U228 ( .A0(n830), .A1(STOP5), .B0(n1357), .B1(STOP6), .Y(n93) );
  INVX1 U229 ( .A(n94), .Y(n762) );
  AOI22X1 U230 ( .A0(n830), .A1(STOP4), .B0(n1336), .B1(STOP5), .Y(n94) );
  INVX1 U231 ( .A(n95), .Y(n763) );
  AOI22X1 U232 ( .A0(n830), .A1(STOP3), .B0(n1384), .B1(STOP4), .Y(n95) );
  INVX1 U233 ( .A(n96), .Y(n764) );
  AOI22X1 U234 ( .A0(n830), .A1(STOP2), .B0(n1356), .B1(STOP3), .Y(n96) );
  INVX1 U235 ( .A(n97), .Y(n765) );
  AOI22X1 U236 ( .A0(n830), .A1(STOP1), .B0(n1355), .B1(STOP2), .Y(n97) );
  INVX1 U237 ( .A(n555), .Y(n1224) );
  AOI22X1 U238 ( .A0(n662), .A1(START5), .B0(n1406), .B1(START6), .Y(n555) );
  INVX1 U239 ( .A(n556), .Y(n1225) );
  AOI22X1 U240 ( .A0(n662), .A1(START4), .B0(n1338), .B1(START5), .Y(n556) );
  INVX1 U241 ( .A(n557), .Y(n1226) );
  AOI22X1 U242 ( .A0(n662), .A1(START3), .B0(n1335), .B1(START4), .Y(n557) );
  INVX1 U243 ( .A(n558), .Y(n1227) );
  AOI22X1 U244 ( .A0(n662), .A1(START2), .B0(n1338), .B1(START3), .Y(n558) );
  INVX1 U245 ( .A(n559), .Y(n1228) );
  AOI22X1 U246 ( .A0(n662), .A1(START1), .B0(n1373), .B1(START2), .Y(n559) );
  INVX1 U247 ( .A(n6), .Y(n674) );
  AOI22X1 U248 ( .A0(DR7[4]), .A1(n649), .B0(DR8[4]), .B1(n1346), .Y(n6) );
  NOR3X1 U249 ( .A(count[0]), .B(count[1]), .C(n1389), .Y(n570) );
  OAI2BB2X1 U250 ( .B0(n646), .B1(n654), .A0N(n1329), .A1N(s_reg[1]), .Y(n756)
         );
  OAI2BB2X1 U251 ( .B0(n646), .B1(n663), .A0N(n1329), .A1N(START7), .Y(n1222)
         );
  OAI2BB2X1 U252 ( .B0(n646), .B1(n651), .A0N(n1329), .A1N(stop3[1]), .Y(n1230) );
  OAI2BB2X1 U253 ( .B0(n646), .B1(n648), .A0N(n1329), .A1N(stop2[1]), .Y(n1233) );
  OAI2BB2X1 U254 ( .B0(n646), .B1(n645), .A0N(n1329), .A1N(stop1[1]), .Y(n1236) );
  OAI2BB2X1 U255 ( .B0(n646), .B1(n672), .A0N(start), .A1N(n1329), .Y(n1302)
         );
  OAI2BB2X1 U256 ( .B0(n646), .B1(n673), .A0N(stop_i), .A1N(n1329), .Y(n1303)
         );
  NAND4X1 U257 ( .A(n2), .B(n3), .C(n4), .D(n5), .Y(out_sel2) );
  NOR3X1 U258 ( .A(out_sel[0]), .B(out_sel[11]), .C(out_sel[10]), .Y(n2) );
  NOR3X1 U259 ( .A(out_sel[12]), .B(out_sel[2]), .C(out_sel[1]), .Y(n3) );
  AOI31X1 U260 ( .A0(n567), .A1(n568), .A2(n569), .B0(n671), .Y(n1239) );
  NOR3X1 U261 ( .A(count[3]), .B(count[6]), .C(count[5]), .Y(n567) );
  NOR3X1 U262 ( .A(count[7]), .B(count[9]), .C(count[8]), .Y(n568) );
  AND3X2 U263 ( .A(n570), .B(count[2]), .C(count[4]), .Y(n569) );
  INVX1 U264 ( .A(n315), .Y(n983) );
  AOI22X1 U265 ( .A0(n1378), .A1(LLL2[12]), .B0(n1320), .B1(LLL1[12]), .Y(n315) );
  INVX1 U266 ( .A(n307), .Y(n975) );
  AOI22X1 U267 ( .A0(n655), .A1(L1[12]), .B0(L2[12]), .B1(n1350), .Y(n307) );
  INVX1 U268 ( .A(n397), .Y(n1065) );
  AOI22X1 U269 ( .A0(n652), .A1(L1[3]), .B0(L2[3]), .B1(n1357), .Y(n397) );
  INVX1 U270 ( .A(n573), .Y(n1242) );
  AOI22X1 U271 ( .A0(n1338), .A1(count[7]), .B0(N183), .B1(n1064), .Y(n573) );
  INVX1 U272 ( .A(n577), .Y(n1246) );
  AOI22X1 U273 ( .A0(n1339), .A1(count[3]), .B0(N179), .B1(n1064), .Y(n577) );
  INVX1 U274 ( .A(n574), .Y(n1243) );
  AOI22X1 U275 ( .A0(n1336), .A1(count[6]), .B0(N182), .B1(n1064), .Y(n574) );
  INVX1 U276 ( .A(n579), .Y(n1248) );
  AOI22X1 U277 ( .A0(n1390), .A1(count[1]), .B0(N177), .B1(n1066), .Y(n579) );
  INVX1 U278 ( .A(n572), .Y(n1241) );
  AOI22X1 U279 ( .A0(n1334), .A1(count[8]), .B0(N184), .B1(n1056), .Y(n572) );
  INVX1 U280 ( .A(n575), .Y(n1244) );
  AOI22X1 U281 ( .A0(n1339), .A1(count[5]), .B0(N181), .B1(n1064), .Y(n575) );
  INVX1 U282 ( .A(n8), .Y(n675) );
  AOI22X1 U283 ( .A0(n1333), .A1(DR7[4]), .B0(n1318), .B1(DR6[4]), .Y(n8) );
  INVX1 U284 ( .A(n9), .Y(n676) );
  AOI22X1 U285 ( .A0(n1337), .A1(DR6[4]), .B0(n1318), .B1(DR5[4]), .Y(n9) );
  INVX1 U286 ( .A(n10), .Y(n677) );
  AOI22X1 U287 ( .A0(n1335), .A1(DR5[4]), .B0(n1316), .B1(DR4[4]), .Y(n10) );
  INVX1 U288 ( .A(n11), .Y(n678) );
  AOI22X1 U289 ( .A0(n1336), .A1(DR4[4]), .B0(n1316), .B1(DR3[4]), .Y(n11) );
  INVX1 U290 ( .A(n12), .Y(n679) );
  AOI22X1 U291 ( .A0(n1335), .A1(DR3[4]), .B0(n1316), .B1(DR2[4]), .Y(n12) );
  INVX1 U292 ( .A(n13), .Y(n680) );
  AOI22X1 U293 ( .A0(n1334), .A1(DR2[4]), .B0(n1317), .B1(DR1[4]), .Y(n13) );
  INVX1 U294 ( .A(n16), .Y(n683) );
  AOI22X1 U295 ( .A0(n1334), .A1(DR7[3]), .B0(n1318), .B1(DR6[3]), .Y(n16) );
  INVX1 U296 ( .A(n17), .Y(n684) );
  AOI22X1 U297 ( .A0(n1406), .A1(DR6[3]), .B0(n1317), .B1(DR5[3]), .Y(n17) );
  INVX1 U298 ( .A(n18), .Y(n685) );
  AOI22X1 U299 ( .A0(n1335), .A1(DR5[3]), .B0(n1318), .B1(DR4[3]), .Y(n18) );
  INVX1 U300 ( .A(n19), .Y(n686) );
  AOI22X1 U301 ( .A0(n1331), .A1(DR4[3]), .B0(n1317), .B1(DR3[3]), .Y(n19) );
  INVX1 U302 ( .A(n20), .Y(n687) );
  AOI22X1 U303 ( .A0(n1405), .A1(DR3[3]), .B0(n1317), .B1(DR2[3]), .Y(n20) );
  INVX1 U304 ( .A(n21), .Y(n688) );
  AOI22X1 U305 ( .A0(n1405), .A1(DR2[3]), .B0(n1318), .B1(DR1[3]), .Y(n21) );
  INVX1 U306 ( .A(n24), .Y(n691) );
  AOI22X1 U307 ( .A0(n1332), .A1(DR7[2]), .B0(n1317), .B1(DR6[2]), .Y(n24) );
  INVX1 U308 ( .A(n25), .Y(n692) );
  AOI22X1 U309 ( .A0(n1331), .A1(DR6[2]), .B0(n1317), .B1(DR5[2]), .Y(n25) );
  INVX1 U310 ( .A(n26), .Y(n693) );
  AOI22X1 U311 ( .A0(n1331), .A1(DR5[2]), .B0(n1317), .B1(DR4[2]), .Y(n26) );
  INVX1 U312 ( .A(n27), .Y(n694) );
  AOI22X1 U313 ( .A0(n1330), .A1(DR4[2]), .B0(n1319), .B1(DR3[2]), .Y(n27) );
  INVX1 U314 ( .A(n28), .Y(n695) );
  AOI22X1 U315 ( .A0(n1333), .A1(DR3[2]), .B0(n1317), .B1(DR2[2]), .Y(n28) );
  INVX1 U316 ( .A(n29), .Y(n696) );
  AOI22X1 U317 ( .A0(n1336), .A1(DR2[2]), .B0(n1317), .B1(DR1[2]), .Y(n29) );
  INVX1 U318 ( .A(n32), .Y(n699) );
  AOI22X1 U319 ( .A0(n1335), .A1(DR7[1]), .B0(n1319), .B1(DR6[1]), .Y(n32) );
  INVX1 U320 ( .A(n33), .Y(n700) );
  AOI22X1 U321 ( .A0(n1332), .A1(DR6[1]), .B0(n1318), .B1(DR5[1]), .Y(n33) );
  INVX1 U322 ( .A(n34), .Y(n701) );
  AOI22X1 U323 ( .A0(n1330), .A1(DR5[1]), .B0(n1318), .B1(DR4[1]), .Y(n34) );
  INVX1 U324 ( .A(n35), .Y(n702) );
  AOI22X1 U325 ( .A0(n1334), .A1(DR4[1]), .B0(n1318), .B1(DR3[1]), .Y(n35) );
  INVX1 U326 ( .A(n36), .Y(n703) );
  AOI22X1 U327 ( .A0(n1335), .A1(DR3[1]), .B0(n1318), .B1(DR2[1]), .Y(n36) );
  INVX1 U328 ( .A(n37), .Y(n704) );
  AOI22X1 U329 ( .A0(n1340), .A1(DR2[1]), .B0(n1318), .B1(DR1[1]), .Y(n37) );
  INVX1 U330 ( .A(n40), .Y(n707) );
  AOI22X1 U331 ( .A0(n1332), .A1(DR7[0]), .B0(n1319), .B1(DR6[0]), .Y(n40) );
  INVX1 U332 ( .A(n41), .Y(n708) );
  AOI22X1 U333 ( .A0(n1336), .A1(DR6[0]), .B0(n1319), .B1(DR5[0]), .Y(n41) );
  INVX1 U334 ( .A(n42), .Y(n709) );
  AOI22X1 U335 ( .A0(n1406), .A1(DR5[0]), .B0(n1319), .B1(DR4[0]), .Y(n42) );
  INVX1 U336 ( .A(n43), .Y(n710) );
  AOI22X1 U337 ( .A0(n1406), .A1(DR4[0]), .B0(n1319), .B1(DR3[0]), .Y(n43) );
  INVX1 U338 ( .A(n44), .Y(n711) );
  AOI22X1 U339 ( .A0(n1340), .A1(DR3[0]), .B0(n1319), .B1(DR2[0]), .Y(n44) );
  INVX1 U340 ( .A(n45), .Y(n712) );
  AOI22X1 U341 ( .A0(n1339), .A1(DR2[0]), .B0(n1319), .B1(DR1[0]), .Y(n45) );
  INVX1 U342 ( .A(n48), .Y(n715) );
  AOI22X1 U343 ( .A0(n1383), .A1(DQ7[4]), .B0(n1319), .B1(DQ6[4]), .Y(n48) );
  INVX1 U344 ( .A(n49), .Y(n716) );
  AOI22X1 U345 ( .A0(n1387), .A1(DQ6[4]), .B0(n1319), .B1(DQ5[4]), .Y(n49) );
  INVX1 U346 ( .A(n50), .Y(n717) );
  AOI22X1 U347 ( .A0(n1331), .A1(DQ5[4]), .B0(n1317), .B1(DQ4[4]), .Y(n50) );
  INVX1 U348 ( .A(n51), .Y(n718) );
  AOI22X1 U349 ( .A0(n1386), .A1(DQ4[4]), .B0(n1327), .B1(DQ3[4]), .Y(n51) );
  INVX1 U350 ( .A(n52), .Y(n719) );
  AOI22X1 U351 ( .A0(n1375), .A1(DQ3[4]), .B0(n1392), .B1(DQ2[4]), .Y(n52) );
  INVX1 U352 ( .A(n53), .Y(n720) );
  AOI22X1 U353 ( .A0(n1382), .A1(DQ2[4]), .B0(n1395), .B1(DQ1[4]), .Y(n53) );
  INVX1 U354 ( .A(n56), .Y(n723) );
  AOI22X1 U355 ( .A0(n1372), .A1(DQ7[3]), .B0(N99), .B1(DQ6[3]), .Y(n56) );
  INVX1 U356 ( .A(n57), .Y(n724) );
  AOI22X1 U357 ( .A0(n1389), .A1(DQ6[3]), .B0(n1394), .B1(DQ5[3]), .Y(n57) );
  INVX1 U358 ( .A(n58), .Y(n725) );
  AOI22X1 U359 ( .A0(n1386), .A1(DQ5[3]), .B0(n1392), .B1(DQ4[3]), .Y(n58) );
  INVX1 U360 ( .A(n59), .Y(n726) );
  AOI22X1 U361 ( .A0(n1375), .A1(DQ4[3]), .B0(n1327), .B1(DQ3[3]), .Y(n59) );
  INVX1 U362 ( .A(n60), .Y(n727) );
  AOI22X1 U363 ( .A0(n1385), .A1(DQ3[3]), .B0(n1396), .B1(DQ2[3]), .Y(n60) );
  INVX1 U364 ( .A(n61), .Y(n728) );
  AOI22X1 U365 ( .A0(n1379), .A1(DQ2[3]), .B0(n1328), .B1(DQ1[3]), .Y(n61) );
  INVX1 U366 ( .A(n64), .Y(n731) );
  AOI22X1 U367 ( .A0(n1372), .A1(DQ7[2]), .B0(n1329), .B1(DQ6[2]), .Y(n64) );
  INVX1 U368 ( .A(n65), .Y(n732) );
  AOI22X1 U369 ( .A0(n1378), .A1(DQ6[2]), .B0(n1328), .B1(DQ5[2]), .Y(n65) );
  INVX1 U370 ( .A(n66), .Y(n733) );
  AOI22X1 U371 ( .A0(n1387), .A1(DQ5[2]), .B0(n1328), .B1(DQ4[2]), .Y(n66) );
  INVX1 U372 ( .A(n67), .Y(n734) );
  AOI22X1 U373 ( .A0(n1335), .A1(DQ4[2]), .B0(n1328), .B1(DQ3[2]), .Y(n67) );
  INVX1 U374 ( .A(n68), .Y(n735) );
  AOI22X1 U375 ( .A0(n1406), .A1(DQ3[2]), .B0(n1329), .B1(DQ2[2]), .Y(n68) );
  INVX1 U376 ( .A(n69), .Y(n736) );
  AOI22X1 U377 ( .A0(n1335), .A1(DQ2[2]), .B0(n1327), .B1(DQ1[2]), .Y(n69) );
  INVX1 U378 ( .A(n72), .Y(n739) );
  AOI22X1 U379 ( .A0(n1339), .A1(DQ7[1]), .B0(n1394), .B1(DQ6[1]), .Y(n72) );
  INVX1 U380 ( .A(n73), .Y(n740) );
  AOI22X1 U381 ( .A0(n1338), .A1(DQ6[1]), .B0(n1328), .B1(DQ5[1]), .Y(n73) );
  INVX1 U382 ( .A(n74), .Y(n741) );
  AOI22X1 U383 ( .A0(n1332), .A1(DQ5[1]), .B0(n1397), .B1(DQ4[1]), .Y(n74) );
  INVX1 U384 ( .A(n75), .Y(n742) );
  AOI22X1 U385 ( .A0(n1333), .A1(DQ4[1]), .B0(n1328), .B1(DQ3[1]), .Y(n75) );
  INVX1 U386 ( .A(n76), .Y(n743) );
  AOI22X1 U387 ( .A0(n1333), .A1(DQ3[1]), .B0(n1329), .B1(DQ2[1]), .Y(n76) );
  INVX1 U388 ( .A(n77), .Y(n744) );
  AOI22X1 U389 ( .A0(n1373), .A1(DQ2[1]), .B0(n1327), .B1(DQ1[1]), .Y(n77) );
  INVX1 U390 ( .A(n80), .Y(n747) );
  AOI22X1 U391 ( .A0(n1385), .A1(DQ7[0]), .B0(n1397), .B1(DQ6[0]), .Y(n80) );
  INVX1 U392 ( .A(n81), .Y(n748) );
  AOI22X1 U393 ( .A0(n1332), .A1(DQ6[0]), .B0(n1328), .B1(DQ5[0]), .Y(n81) );
  INVX1 U394 ( .A(n82), .Y(n749) );
  AOI22X1 U395 ( .A0(n1330), .A1(DQ5[0]), .B0(n1399), .B1(DQ4[0]), .Y(n82) );
  INVX1 U396 ( .A(n83), .Y(n750) );
  AOI22X1 U397 ( .A0(n1332), .A1(DQ4[0]), .B0(n1327), .B1(DQ3[0]), .Y(n83) );
  INVX1 U398 ( .A(n84), .Y(n751) );
  AOI22X1 U399 ( .A0(n1338), .A1(DQ3[0]), .B0(n1393), .B1(DQ2[0]), .Y(n84) );
  INVX1 U400 ( .A(n85), .Y(n752) );
  AOI22X1 U401 ( .A0(n1341), .A1(DQ2[0]), .B0(n1326), .B1(DQ1[0]), .Y(n85) );
  INVX1 U402 ( .A(n100), .Y(n768) );
  AOI22X1 U403 ( .A0(n830), .A1(R6[12]), .B0(n1365), .B1(R7[12]), .Y(n100) );
  INVX1 U404 ( .A(n101), .Y(n769) );
  AOI22X1 U405 ( .A0(n830), .A1(R5[12]), .B0(n1366), .B1(R6[12]), .Y(n101) );
  INVX1 U406 ( .A(n102), .Y(n770) );
  AOI22X1 U407 ( .A0(n830), .A1(R4[12]), .B0(n1364), .B1(R5[12]), .Y(n102) );
  INVX1 U408 ( .A(n103), .Y(n771) );
  AOI22X1 U409 ( .A0(n838), .A1(R3[12]), .B0(n1344), .B1(R4[12]), .Y(n103) );
  INVX1 U410 ( .A(n104), .Y(n772) );
  AOI22X1 U411 ( .A0(n838), .A1(R2[12]), .B0(n1348), .B1(R3[12]), .Y(n104) );
  INVX1 U412 ( .A(n105), .Y(n773) );
  AOI22X1 U413 ( .A0(n838), .A1(R1[12]), .B0(n1349), .B1(R2[12]), .Y(n105) );
  INVX1 U414 ( .A(n108), .Y(n776) );
  AOI22X1 U415 ( .A0(n838), .A1(R6[11]), .B0(n1345), .B1(R7[11]), .Y(n108) );
  INVX1 U416 ( .A(n109), .Y(n777) );
  AOI22X1 U417 ( .A0(n838), .A1(R5[11]), .B0(n1351), .B1(R6[11]), .Y(n109) );
  INVX1 U418 ( .A(n110), .Y(n778) );
  AOI22X1 U419 ( .A0(n838), .A1(R4[11]), .B0(n1361), .B1(R5[11]), .Y(n110) );
  INVX1 U420 ( .A(n111), .Y(n779) );
  AOI22X1 U421 ( .A0(n838), .A1(R3[11]), .B0(n1390), .B1(R4[11]), .Y(n111) );
  INVX1 U422 ( .A(n112), .Y(n780) );
  AOI22X1 U423 ( .A0(n838), .A1(R2[11]), .B0(n1347), .B1(R3[11]), .Y(n112) );
  INVX1 U424 ( .A(n113), .Y(n781) );
  AOI22X1 U425 ( .A0(n838), .A1(R1[11]), .B0(n1377), .B1(R2[11]), .Y(n113) );
  INVX1 U426 ( .A(n116), .Y(n784) );
  AOI22X1 U427 ( .A0(n846), .A1(R6[10]), .B0(n1343), .B1(R7[10]), .Y(n116) );
  INVX1 U428 ( .A(n117), .Y(n785) );
  AOI22X1 U429 ( .A0(n846), .A1(R5[10]), .B0(n1363), .B1(R6[10]), .Y(n117) );
  INVX1 U430 ( .A(n118), .Y(n786) );
  AOI22X1 U431 ( .A0(n846), .A1(R4[10]), .B0(n1364), .B1(R5[10]), .Y(n118) );
  INVX1 U432 ( .A(n119), .Y(n787) );
  AOI22X1 U433 ( .A0(n846), .A1(R3[10]), .B0(n1365), .B1(R4[10]), .Y(n119) );
  INVX1 U434 ( .A(n120), .Y(n788) );
  AOI22X1 U435 ( .A0(n846), .A1(R2[10]), .B0(n1346), .B1(R3[10]), .Y(n120) );
  INVX1 U436 ( .A(n121), .Y(n789) );
  AOI22X1 U437 ( .A0(n846), .A1(R1[10]), .B0(n1363), .B1(R2[10]), .Y(n121) );
  INVX1 U438 ( .A(n124), .Y(n792) );
  AOI22X1 U439 ( .A0(n846), .A1(R6[9]), .B0(n1346), .B1(R7[9]), .Y(n124) );
  INVX1 U440 ( .A(n125), .Y(n793) );
  AOI22X1 U441 ( .A0(n846), .A1(R5[9]), .B0(n1365), .B1(R6[9]), .Y(n125) );
  INVX1 U442 ( .A(n126), .Y(n794) );
  AOI22X1 U443 ( .A0(n986), .A1(R4[9]), .B0(n1364), .B1(R5[9]), .Y(n126) );
  INVX1 U444 ( .A(n127), .Y(n795) );
  AOI22X1 U445 ( .A0(n986), .A1(R3[9]), .B0(n1353), .B1(R4[9]), .Y(n127) );
  INVX1 U446 ( .A(n128), .Y(n796) );
  AOI22X1 U447 ( .A0(n986), .A1(R2[9]), .B0(n1359), .B1(R3[9]), .Y(n128) );
  INVX1 U448 ( .A(n129), .Y(n797) );
  AOI22X1 U449 ( .A0(n986), .A1(R1[9]), .B0(n1356), .B1(R2[9]), .Y(n129) );
  INVX1 U450 ( .A(n132), .Y(n800) );
  AOI22X1 U451 ( .A0(n986), .A1(R6[8]), .B0(n1354), .B1(R7[8]), .Y(n132) );
  INVX1 U452 ( .A(n133), .Y(n801) );
  AOI22X1 U453 ( .A0(n986), .A1(R5[8]), .B0(n1356), .B1(R6[8]), .Y(n133) );
  INVX1 U454 ( .A(n134), .Y(n802) );
  AOI22X1 U455 ( .A0(n986), .A1(R4[8]), .B0(n1352), .B1(R5[8]), .Y(n134) );
  INVX1 U456 ( .A(n135), .Y(n803) );
  AOI22X1 U457 ( .A0(n986), .A1(R3[8]), .B0(n1366), .B1(R4[8]), .Y(n135) );
  INVX1 U458 ( .A(n136), .Y(n804) );
  AOI22X1 U459 ( .A0(n986), .A1(R2[8]), .B0(n1368), .B1(R3[8]), .Y(n136) );
  INVX1 U460 ( .A(n137), .Y(n805) );
  AOI22X1 U461 ( .A0(n994), .A1(R1[8]), .B0(n1354), .B1(R2[8]), .Y(n137) );
  INVX1 U462 ( .A(n140), .Y(n808) );
  AOI22X1 U463 ( .A0(n994), .A1(R6[7]), .B0(n1350), .B1(R7[7]), .Y(n140) );
  INVX1 U464 ( .A(n141), .Y(n809) );
  AOI22X1 U465 ( .A0(n994), .A1(R5[7]), .B0(n1350), .B1(R6[7]), .Y(n141) );
  INVX1 U466 ( .A(n142), .Y(n810) );
  AOI22X1 U467 ( .A0(n994), .A1(R4[7]), .B0(n1400), .B1(R5[7]), .Y(n142) );
  INVX1 U468 ( .A(n143), .Y(n811) );
  AOI22X1 U469 ( .A0(n994), .A1(R3[7]), .B0(n1337), .B1(R4[7]), .Y(n143) );
  INVX1 U470 ( .A(n144), .Y(n812) );
  AOI22X1 U471 ( .A0(n994), .A1(R2[7]), .B0(n1343), .B1(R3[7]), .Y(n144) );
  INVX1 U472 ( .A(n145), .Y(n813) );
  AOI22X1 U473 ( .A0(n994), .A1(R1[7]), .B0(n1370), .B1(R2[7]), .Y(n145) );
  INVX1 U474 ( .A(n148), .Y(n816) );
  AOI22X1 U475 ( .A0(n994), .A1(R6[6]), .B0(n1402), .B1(R7[6]), .Y(n148) );
  INVX1 U476 ( .A(n149), .Y(n817) );
  AOI22X1 U477 ( .A0(n996), .A1(R5[6]), .B0(n1405), .B1(R6[6]), .Y(n149) );
  INVX1 U478 ( .A(n150), .Y(n818) );
  AOI22X1 U479 ( .A0(n996), .A1(R4[6]), .B0(n1408), .B1(R5[6]), .Y(n150) );
  INVX1 U480 ( .A(n151), .Y(n819) );
  AOI22X1 U481 ( .A0(n996), .A1(R3[6]), .B0(n1380), .B1(R4[6]), .Y(n151) );
  INVX1 U482 ( .A(n152), .Y(n820) );
  AOI22X1 U483 ( .A0(n996), .A1(R2[6]), .B0(n1338), .B1(R3[6]), .Y(n152) );
  INVX1 U484 ( .A(n153), .Y(n821) );
  AOI22X1 U485 ( .A0(n996), .A1(R1[6]), .B0(n1370), .B1(R2[6]), .Y(n153) );
  INVX1 U486 ( .A(n156), .Y(n824) );
  AOI22X1 U487 ( .A0(n996), .A1(R6[5]), .B0(n1342), .B1(R7[5]), .Y(n156) );
  INVX1 U488 ( .A(n157), .Y(n825) );
  AOI22X1 U489 ( .A0(n996), .A1(R5[5]), .B0(n1345), .B1(R6[5]), .Y(n157) );
  INVX1 U490 ( .A(n158), .Y(n826) );
  AOI22X1 U491 ( .A0(n996), .A1(R4[5]), .B0(n1406), .B1(R5[5]), .Y(n158) );
  INVX1 U492 ( .A(n159), .Y(n827) );
  AOI22X1 U493 ( .A0(n996), .A1(R3[5]), .B0(n1360), .B1(R4[5]), .Y(n159) );
  INVX1 U494 ( .A(n160), .Y(n828) );
  AOI22X1 U495 ( .A0(n1004), .A1(R2[5]), .B0(n1403), .B1(R3[5]), .Y(n160) );
  INVX1 U496 ( .A(n161), .Y(n829) );
  AOI22X1 U497 ( .A0(n1004), .A1(R1[5]), .B0(n1385), .B1(R2[5]), .Y(n161) );
  INVX1 U498 ( .A(n164), .Y(n832) );
  AOI22X1 U499 ( .A0(n1004), .A1(R6[4]), .B0(n1345), .B1(R7[4]), .Y(n164) );
  INVX1 U500 ( .A(n165), .Y(n833) );
  AOI22X1 U501 ( .A0(n1004), .A1(R5[4]), .B0(n1400), .B1(R6[4]), .Y(n165) );
  INVX1 U502 ( .A(n166), .Y(n834) );
  AOI22X1 U503 ( .A0(n1004), .A1(R4[4]), .B0(n1402), .B1(R5[4]), .Y(n166) );
  INVX1 U504 ( .A(n167), .Y(n835) );
  AOI22X1 U505 ( .A0(n1006), .A1(R3[4]), .B0(n1406), .B1(R4[4]), .Y(n167) );
  INVX1 U506 ( .A(n168), .Y(n836) );
  AOI22X1 U507 ( .A0(n1014), .A1(R2[4]), .B0(n1341), .B1(R3[4]), .Y(n168) );
  INVX1 U508 ( .A(n169), .Y(n837) );
  AOI22X1 U509 ( .A0(n1016), .A1(R1[4]), .B0(n1370), .B1(R2[4]), .Y(n169) );
  INVX1 U510 ( .A(n172), .Y(n840) );
  AOI22X1 U511 ( .A0(n1006), .A1(R6[3]), .B0(n1384), .B1(R7[3]), .Y(n172) );
  INVX1 U512 ( .A(n173), .Y(n841) );
  AOI22X1 U513 ( .A0(n1024), .A1(R5[3]), .B0(n1338), .B1(R6[3]), .Y(n173) );
  INVX1 U514 ( .A(n174), .Y(n842) );
  AOI22X1 U515 ( .A0(n1014), .A1(R4[3]), .B0(n1373), .B1(R5[3]), .Y(n174) );
  INVX1 U516 ( .A(n175), .Y(n843) );
  AOI22X1 U517 ( .A0(n1016), .A1(R3[3]), .B0(n1353), .B1(R4[3]), .Y(n175) );
  INVX1 U518 ( .A(n176), .Y(n844) );
  AOI22X1 U519 ( .A0(n1026), .A1(R2[3]), .B0(n1379), .B1(R3[3]), .Y(n176) );
  INVX1 U520 ( .A(n177), .Y(n845) );
  AOI22X1 U521 ( .A0(n1026), .A1(R1[3]), .B0(n1375), .B1(R2[3]), .Y(n177) );
  INVX1 U522 ( .A(n180), .Y(n848) );
  AOI22X1 U523 ( .A0(n1034), .A1(R6[2]), .B0(n1355), .B1(R7[2]), .Y(n180) );
  INVX1 U524 ( .A(n181), .Y(n849) );
  AOI22X1 U525 ( .A0(n1024), .A1(R5[2]), .B0(n1360), .B1(R6[2]), .Y(n181) );
  INVX1 U526 ( .A(n182), .Y(n850) );
  AOI22X1 U527 ( .A0(n1034), .A1(R4[2]), .B0(n1367), .B1(R5[2]), .Y(n182) );
  INVX1 U528 ( .A(n183), .Y(n851) );
  AOI22X1 U529 ( .A0(n1026), .A1(R3[2]), .B0(n1358), .B1(R4[2]), .Y(n183) );
  INVX1 U530 ( .A(n184), .Y(n852) );
  AOI22X1 U531 ( .A0(n1006), .A1(R2[2]), .B0(n1357), .B1(R3[2]), .Y(n184) );
  INVX1 U532 ( .A(n185), .Y(n853) );
  AOI22X1 U533 ( .A0(n1034), .A1(R1[2]), .B0(n1375), .B1(R2[2]), .Y(n185) );
  INVX1 U534 ( .A(n188), .Y(n856) );
  AOI22X1 U535 ( .A0(n1034), .A1(R6[1]), .B0(n1375), .B1(R7[1]), .Y(n188) );
  INVX1 U536 ( .A(n189), .Y(n857) );
  AOI22X1 U537 ( .A0(n1034), .A1(R5[1]), .B0(n1369), .B1(R6[1]), .Y(n189) );
  INVX1 U538 ( .A(n190), .Y(n858) );
  AOI22X1 U539 ( .A0(n1024), .A1(R4[1]), .B0(n1362), .B1(R5[1]), .Y(n190) );
  INVX1 U540 ( .A(n191), .Y(n859) );
  AOI22X1 U541 ( .A0(n1026), .A1(R3[1]), .B0(n1371), .B1(R4[1]), .Y(n191) );
  INVX1 U542 ( .A(n192), .Y(n860) );
  AOI22X1 U543 ( .A0(n1024), .A1(R2[1]), .B0(n1339), .B1(R3[1]), .Y(n192) );
  INVX1 U544 ( .A(n193), .Y(n861) );
  AOI22X1 U545 ( .A0(n1034), .A1(R1[1]), .B0(n1348), .B1(R2[1]), .Y(n193) );
  INVX1 U546 ( .A(n196), .Y(n864) );
  AOI22X1 U547 ( .A0(n1026), .A1(R6[0]), .B0(n1361), .B1(R7[0]), .Y(n196) );
  INVX1 U548 ( .A(n197), .Y(n865) );
  AOI22X1 U549 ( .A0(n1026), .A1(R5[0]), .B0(n1358), .B1(R6[0]), .Y(n197) );
  INVX1 U550 ( .A(n198), .Y(n866) );
  AOI22X1 U551 ( .A0(n1016), .A1(R4[0]), .B0(n1341), .B1(R5[0]), .Y(n198) );
  INVX1 U552 ( .A(n199), .Y(n867) );
  AOI22X1 U553 ( .A0(n1026), .A1(R3[0]), .B0(n1336), .B1(R4[0]), .Y(n199) );
  INVX1 U554 ( .A(n200), .Y(n868) );
  AOI22X1 U555 ( .A0(n1016), .A1(R2[0]), .B0(n1346), .B1(R3[0]), .Y(n200) );
  INVX1 U556 ( .A(n201), .Y(n869) );
  AOI22X1 U557 ( .A0(n1026), .A1(R1[0]), .B0(n1346), .B1(R2[0]), .Y(n201) );
  INVX1 U558 ( .A(n204), .Y(n872) );
  AOI22X1 U559 ( .A0(n1016), .A1(Q6[12]), .B0(n1361), .B1(Q7[12]), .Y(n204) );
  INVX1 U560 ( .A(n205), .Y(n873) );
  AOI22X1 U561 ( .A0(n1016), .A1(Q5[12]), .B0(n1342), .B1(Q6[12]), .Y(n205) );
  INVX1 U562 ( .A(n206), .Y(n874) );
  AOI22X1 U563 ( .A0(n1024), .A1(Q4[12]), .B0(n1380), .B1(Q5[12]), .Y(n206) );
  INVX1 U564 ( .A(n207), .Y(n875) );
  AOI22X1 U565 ( .A0(n1016), .A1(Q3[12]), .B0(n1389), .B1(Q4[12]), .Y(n207) );
  INVX1 U566 ( .A(n208), .Y(n876) );
  AOI22X1 U567 ( .A0(n1024), .A1(Q2[12]), .B0(n1363), .B1(Q3[12]), .Y(n208) );
  INVX1 U568 ( .A(n209), .Y(n877) );
  AOI22X1 U569 ( .A0(n1024), .A1(Q1[12]), .B0(n1361), .B1(Q2[12]), .Y(n209) );
  INVX1 U570 ( .A(n212), .Y(n880) );
  AOI22X1 U571 ( .A0(n1024), .A1(Q6[11]), .B0(n1342), .B1(Q7[11]), .Y(n212) );
  INVX1 U572 ( .A(n213), .Y(n881) );
  AOI22X1 U573 ( .A0(n1014), .A1(Q5[11]), .B0(n1408), .B1(Q6[11]), .Y(n213) );
  INVX1 U574 ( .A(n214), .Y(n882) );
  AOI22X1 U575 ( .A0(n1014), .A1(Q4[11]), .B0(n1361), .B1(Q5[11]), .Y(n214) );
  INVX1 U576 ( .A(n215), .Y(n883) );
  AOI22X1 U577 ( .A0(n1016), .A1(Q3[11]), .B0(n1349), .B1(Q4[11]), .Y(n215) );
  INVX1 U578 ( .A(n216), .Y(n884) );
  AOI22X1 U579 ( .A0(n1016), .A1(Q2[11]), .B0(n1372), .B1(Q3[11]), .Y(n216) );
  INVX1 U580 ( .A(n217), .Y(n885) );
  AOI22X1 U581 ( .A0(n1006), .A1(Q1[11]), .B0(n1348), .B1(Q2[11]), .Y(n217) );
  INVX1 U582 ( .A(n220), .Y(n888) );
  AOI22X1 U583 ( .A0(n1006), .A1(Q6[10]), .B0(n1349), .B1(Q7[10]), .Y(n220) );
  INVX1 U584 ( .A(n221), .Y(n889) );
  AOI22X1 U585 ( .A0(n1014), .A1(Q5[10]), .B0(n1383), .B1(Q6[10]), .Y(n221) );
  INVX1 U586 ( .A(n222), .Y(n890) );
  AOI22X1 U587 ( .A0(n1014), .A1(Q4[10]), .B0(n1368), .B1(Q5[10]), .Y(n222) );
  INVX1 U588 ( .A(n223), .Y(n891) );
  AOI22X1 U589 ( .A0(n1006), .A1(Q3[10]), .B0(n1341), .B1(Q4[10]), .Y(n223) );
  INVX1 U590 ( .A(n224), .Y(n892) );
  AOI22X1 U591 ( .A0(n1014), .A1(Q2[10]), .B0(n1389), .B1(Q3[10]), .Y(n224) );
  INVX1 U592 ( .A(n225), .Y(n893) );
  AOI22X1 U593 ( .A0(n1014), .A1(Q1[10]), .B0(n1344), .B1(Q2[10]), .Y(n225) );
  INVX1 U594 ( .A(n228), .Y(n896) );
  AOI22X1 U595 ( .A0(n1006), .A1(Q6[9]), .B0(n1332), .B1(Q7[9]), .Y(n228) );
  INVX1 U596 ( .A(n229), .Y(n897) );
  AOI22X1 U597 ( .A0(n1004), .A1(Q5[9]), .B0(n1367), .B1(Q6[9]), .Y(n229) );
  INVX1 U598 ( .A(n230), .Y(n898) );
  AOI22X1 U599 ( .A0(n1004), .A1(Q4[9]), .B0(n1362), .B1(Q5[9]), .Y(n230) );
  INVX1 U600 ( .A(n231), .Y(n899) );
  AOI22X1 U601 ( .A0(n1006), .A1(Q3[9]), .B0(n1376), .B1(Q4[9]), .Y(n231) );
  INVX1 U602 ( .A(n232), .Y(n900) );
  AOI22X1 U603 ( .A0(n1006), .A1(Q2[9]), .B0(n1366), .B1(Q3[9]), .Y(n232) );
  INVX1 U604 ( .A(n233), .Y(n901) );
  AOI22X1 U605 ( .A0(n1014), .A1(Q1[9]), .B0(n1347), .B1(Q2[9]), .Y(n233) );
  INVX1 U606 ( .A(n236), .Y(n904) );
  AOI22X1 U607 ( .A0(n662), .A1(Q6[8]), .B0(n1369), .B1(Q7[8]), .Y(n236) );
  INVX1 U608 ( .A(n237), .Y(n905) );
  AOI22X1 U609 ( .A0(n662), .A1(Q5[8]), .B0(n1343), .B1(Q6[8]), .Y(n237) );
  INVX1 U610 ( .A(n238), .Y(n906) );
  AOI22X1 U611 ( .A0(n662), .A1(Q4[8]), .B0(n1345), .B1(Q5[8]), .Y(n238) );
  INVX1 U612 ( .A(n239), .Y(n907) );
  AOI22X1 U613 ( .A0(n661), .A1(Q3[8]), .B0(n1351), .B1(Q4[8]), .Y(n239) );
  INVX1 U614 ( .A(n240), .Y(n908) );
  AOI22X1 U615 ( .A0(n661), .A1(Q2[8]), .B0(n1350), .B1(Q3[8]), .Y(n240) );
  INVX1 U616 ( .A(n241), .Y(n909) );
  AOI22X1 U617 ( .A0(n661), .A1(Q1[8]), .B0(n1338), .B1(Q2[8]), .Y(n241) );
  INVX1 U618 ( .A(n244), .Y(n912) );
  AOI22X1 U619 ( .A0(n661), .A1(Q6[7]), .B0(n1348), .B1(Q7[7]), .Y(n244) );
  INVX1 U620 ( .A(n245), .Y(n913) );
  AOI22X1 U621 ( .A0(n661), .A1(Q5[7]), .B0(n1402), .B1(Q6[7]), .Y(n245) );
  INVX1 U622 ( .A(n246), .Y(n914) );
  AOI22X1 U623 ( .A0(n661), .A1(Q4[7]), .B0(n1382), .B1(Q5[7]), .Y(n246) );
  INVX1 U624 ( .A(n247), .Y(n915) );
  AOI22X1 U625 ( .A0(n661), .A1(Q3[7]), .B0(n1341), .B1(Q4[7]), .Y(n247) );
  INVX1 U626 ( .A(n248), .Y(n916) );
  AOI22X1 U627 ( .A0(n661), .A1(Q2[7]), .B0(n1379), .B1(Q3[7]), .Y(n248) );
  INVX1 U628 ( .A(n249), .Y(n917) );
  AOI22X1 U629 ( .A0(n661), .A1(Q1[7]), .B0(n1339), .B1(Q2[7]), .Y(n249) );
  INVX1 U630 ( .A(n252), .Y(n920) );
  AOI22X1 U631 ( .A0(n660), .A1(Q6[6]), .B0(n1340), .B1(Q7[6]), .Y(n252) );
  INVX1 U632 ( .A(n253), .Y(n921) );
  AOI22X1 U633 ( .A0(n660), .A1(Q5[6]), .B0(n1400), .B1(Q6[6]), .Y(n253) );
  INVX1 U634 ( .A(n254), .Y(n922) );
  AOI22X1 U635 ( .A0(n660), .A1(Q4[6]), .B0(n1358), .B1(Q5[6]), .Y(n254) );
  INVX1 U636 ( .A(n255), .Y(n923) );
  AOI22X1 U637 ( .A0(n660), .A1(Q3[6]), .B0(n1351), .B1(Q4[6]), .Y(n255) );
  INVX1 U638 ( .A(n256), .Y(n924) );
  AOI22X1 U639 ( .A0(n660), .A1(Q2[6]), .B0(n1357), .B1(Q3[6]), .Y(n256) );
  INVX1 U640 ( .A(n257), .Y(n925) );
  AOI22X1 U641 ( .A0(n660), .A1(Q1[6]), .B0(n1344), .B1(Q2[6]), .Y(n257) );
  INVX1 U642 ( .A(n260), .Y(n928) );
  AOI22X1 U643 ( .A0(n660), .A1(Q6[5]), .B0(n1339), .B1(Q7[5]), .Y(n260) );
  INVX1 U644 ( .A(n261), .Y(n929) );
  AOI22X1 U645 ( .A0(n660), .A1(Q5[5]), .B0(n1368), .B1(Q6[5]), .Y(n261) );
  INVX1 U646 ( .A(n262), .Y(n930) );
  AOI22X1 U647 ( .A0(n659), .A1(Q4[5]), .B0(n1372), .B1(Q5[5]), .Y(n262) );
  INVX1 U648 ( .A(n263), .Y(n931) );
  AOI22X1 U649 ( .A0(n659), .A1(Q3[5]), .B0(n1381), .B1(Q4[5]), .Y(n263) );
  INVX1 U650 ( .A(n264), .Y(n932) );
  AOI22X1 U651 ( .A0(n659), .A1(Q2[5]), .B0(n1345), .B1(Q3[5]), .Y(n264) );
  INVX1 U652 ( .A(n265), .Y(n933) );
  AOI22X1 U653 ( .A0(n659), .A1(Q1[5]), .B0(n1343), .B1(Q2[5]), .Y(n265) );
  INVX1 U654 ( .A(n268), .Y(n936) );
  AOI22X1 U655 ( .A0(n659), .A1(Q6[4]), .B0(n1347), .B1(Q7[4]), .Y(n268) );
  INVX1 U656 ( .A(n269), .Y(n937) );
  AOI22X1 U657 ( .A0(n659), .A1(Q5[4]), .B0(n1355), .B1(Q6[4]), .Y(n269) );
  INVX1 U658 ( .A(n270), .Y(n938) );
  AOI22X1 U659 ( .A0(n659), .A1(Q4[4]), .B0(n1344), .B1(Q5[4]), .Y(n270) );
  INVX1 U660 ( .A(n271), .Y(n939) );
  AOI22X1 U661 ( .A0(n659), .A1(Q3[4]), .B0(n1337), .B1(Q4[4]), .Y(n271) );
  INVX1 U662 ( .A(n272), .Y(n940) );
  AOI22X1 U663 ( .A0(n659), .A1(Q2[4]), .B0(n1356), .B1(Q3[4]), .Y(n272) );
  INVX1 U664 ( .A(n273), .Y(n941) );
  AOI22X1 U665 ( .A0(n658), .A1(Q1[4]), .B0(n1373), .B1(Q2[4]), .Y(n273) );
  INVX1 U666 ( .A(n276), .Y(n944) );
  AOI22X1 U667 ( .A0(n658), .A1(Q6[3]), .B0(n1381), .B1(Q7[3]), .Y(n276) );
  INVX1 U668 ( .A(n277), .Y(n945) );
  AOI22X1 U669 ( .A0(n658), .A1(Q5[3]), .B0(n1383), .B1(Q6[3]), .Y(n277) );
  INVX1 U670 ( .A(n278), .Y(n946) );
  AOI22X1 U671 ( .A0(n658), .A1(Q4[3]), .B0(n1378), .B1(Q5[3]), .Y(n278) );
  INVX1 U672 ( .A(n279), .Y(n947) );
  AOI22X1 U673 ( .A0(n658), .A1(Q3[3]), .B0(n1345), .B1(Q4[3]), .Y(n279) );
  INVX1 U674 ( .A(n280), .Y(n948) );
  AOI22X1 U675 ( .A0(n658), .A1(Q2[3]), .B0(n1374), .B1(Q3[3]), .Y(n280) );
  INVX1 U676 ( .A(n281), .Y(n949) );
  AOI22X1 U677 ( .A0(n658), .A1(Q1[3]), .B0(n1377), .B1(Q2[3]), .Y(n281) );
  INVX1 U678 ( .A(n284), .Y(n952) );
  AOI22X1 U679 ( .A0(n658), .A1(Q6[2]), .B0(n1354), .B1(Q7[2]), .Y(n284) );
  INVX1 U680 ( .A(n285), .Y(n953) );
  AOI22X1 U681 ( .A0(n657), .A1(Q5[2]), .B0(n1337), .B1(Q6[2]), .Y(n285) );
  INVX1 U682 ( .A(n286), .Y(n954) );
  AOI22X1 U683 ( .A0(n657), .A1(Q4[2]), .B0(n1344), .B1(Q5[2]), .Y(n286) );
  INVX1 U684 ( .A(n287), .Y(n955) );
  AOI22X1 U685 ( .A0(n657), .A1(Q3[2]), .B0(n1400), .B1(Q4[2]), .Y(n287) );
  INVX1 U686 ( .A(n288), .Y(n956) );
  AOI22X1 U687 ( .A0(n657), .A1(Q2[2]), .B0(n1343), .B1(Q3[2]), .Y(n288) );
  INVX1 U688 ( .A(n289), .Y(n957) );
  AOI22X1 U689 ( .A0(n657), .A1(Q1[2]), .B0(n1364), .B1(Q2[2]), .Y(n289) );
  INVX1 U690 ( .A(n292), .Y(n960) );
  AOI22X1 U691 ( .A0(n657), .A1(Q6[1]), .B0(n1341), .B1(Q7[1]), .Y(n292) );
  INVX1 U692 ( .A(n293), .Y(n961) );
  AOI22X1 U693 ( .A0(n657), .A1(Q5[1]), .B0(n1351), .B1(Q6[1]), .Y(n293) );
  INVX1 U694 ( .A(n294), .Y(n962) );
  AOI22X1 U695 ( .A0(n657), .A1(Q4[1]), .B0(n1349), .B1(Q5[1]), .Y(n294) );
  INVX1 U696 ( .A(n295), .Y(n963) );
  AOI22X1 U697 ( .A0(n657), .A1(Q3[1]), .B0(n1369), .B1(Q4[1]), .Y(n295) );
  INVX1 U698 ( .A(n296), .Y(n964) );
  AOI22X1 U699 ( .A0(n656), .A1(Q2[1]), .B0(n1371), .B1(Q3[1]), .Y(n296) );
  INVX1 U700 ( .A(n297), .Y(n965) );
  AOI22X1 U701 ( .A0(n656), .A1(Q1[1]), .B0(n1347), .B1(Q2[1]), .Y(n297) );
  INVX1 U702 ( .A(n300), .Y(n968) );
  AOI22X1 U703 ( .A0(n656), .A1(Q6[0]), .B0(n1330), .B1(Q7[0]), .Y(n300) );
  INVX1 U704 ( .A(n301), .Y(n969) );
  AOI22X1 U705 ( .A0(n656), .A1(Q5[0]), .B0(n1387), .B1(Q6[0]), .Y(n301) );
  INVX1 U706 ( .A(n302), .Y(n970) );
  AOI22X1 U707 ( .A0(n656), .A1(Q4[0]), .B0(n1346), .B1(Q5[0]), .Y(n302) );
  INVX1 U708 ( .A(n303), .Y(n971) );
  AOI22X1 U709 ( .A0(n656), .A1(Q3[0]), .B0(n1400), .B1(Q4[0]), .Y(n303) );
  INVX1 U710 ( .A(n304), .Y(n972) );
  AOI22X1 U711 ( .A0(n656), .A1(Q2[0]), .B0(n1381), .B1(Q3[0]), .Y(n304) );
  INVX1 U712 ( .A(n305), .Y(n973) );
  AOI22X1 U713 ( .A0(n656), .A1(Q1[0]), .B0(n1366), .B1(Q2[0]), .Y(n305) );
  INVX1 U714 ( .A(n310), .Y(n978) );
  AOI22X1 U715 ( .A0(n1361), .A1(LLL7[12]), .B0(n1321), .B1(LLL6[12]), .Y(n310) );
  INVX1 U716 ( .A(n311), .Y(n979) );
  AOI22X1 U717 ( .A0(n1341), .A1(LLL6[12]), .B0(n1321), .B1(LLL5[12]), .Y(n311) );
  INVX1 U718 ( .A(n312), .Y(n980) );
  AOI22X1 U719 ( .A0(n1374), .A1(LLL5[12]), .B0(n1320), .B1(LLL4[12]), .Y(n312) );
  INVX1 U720 ( .A(n313), .Y(n981) );
  AOI22X1 U721 ( .A0(n1390), .A1(LLL4[12]), .B0(n1320), .B1(LLL3[12]), .Y(n313) );
  INVX1 U722 ( .A(n314), .Y(n982) );
  AOI22X1 U723 ( .A0(n1408), .A1(LLL3[12]), .B0(n1326), .B1(LLL2[12]), .Y(n314) );
  INVX1 U724 ( .A(n320), .Y(n988) );
  AOI22X1 U725 ( .A0(n1334), .A1(LLL7[11]), .B0(n1320), .B1(LLL6[11]), .Y(n320) );
  INVX1 U726 ( .A(n321), .Y(n989) );
  AOI22X1 U727 ( .A0(n1408), .A1(LLL6[11]), .B0(n1320), .B1(LLL5[11]), .Y(n321) );
  INVX1 U728 ( .A(n322), .Y(n990) );
  AOI22X1 U729 ( .A0(n1377), .A1(LLL5[11]), .B0(n1320), .B1(LLL4[11]), .Y(n322) );
  INVX1 U730 ( .A(n323), .Y(n991) );
  AOI22X1 U731 ( .A0(n1373), .A1(LLL4[11]), .B0(n1320), .B1(LLL3[11]), .Y(n323) );
  INVX1 U732 ( .A(n324), .Y(n992) );
  AOI22X1 U733 ( .A0(n1365), .A1(LLL3[11]), .B0(n1320), .B1(LLL2[11]), .Y(n324) );
  INVX1 U734 ( .A(n330), .Y(n998) );
  AOI22X1 U735 ( .A0(n1368), .A1(LLL7[10]), .B0(n1321), .B1(LLL6[10]), .Y(n330) );
  INVX1 U736 ( .A(n331), .Y(n999) );
  AOI22X1 U737 ( .A0(n1371), .A1(LLL6[10]), .B0(n1321), .B1(LLL5[10]), .Y(n331) );
  INVX1 U738 ( .A(n332), .Y(n1000) );
  AOI22X1 U739 ( .A0(n1351), .A1(LLL5[10]), .B0(n1321), .B1(LLL4[10]), .Y(n332) );
  INVX1 U740 ( .A(n333), .Y(n1001) );
  AOI22X1 U741 ( .A0(n1350), .A1(LLL4[10]), .B0(n1321), .B1(LLL3[10]), .Y(n333) );
  INVX1 U742 ( .A(n334), .Y(n1002) );
  AOI22X1 U743 ( .A0(n1330), .A1(LLL3[10]), .B0(n1321), .B1(LLL2[10]), .Y(n334) );
  INVX1 U744 ( .A(n340), .Y(n1008) );
  AOI22X1 U745 ( .A0(n1369), .A1(LLL7[9]), .B0(n1321), .B1(LLL6[9]), .Y(n340)
         );
  INVX1 U746 ( .A(n341), .Y(n1009) );
  AOI22X1 U747 ( .A0(n1358), .A1(LLL6[9]), .B0(n1321), .B1(LLL5[9]), .Y(n341)
         );
  INVX1 U748 ( .A(n342), .Y(n1010) );
  AOI22X1 U749 ( .A0(n1334), .A1(LLL5[9]), .B0(n1322), .B1(LLL4[9]), .Y(n342)
         );
  INVX1 U750 ( .A(n343), .Y(n1011) );
  AOI22X1 U751 ( .A0(n1371), .A1(LLL4[9]), .B0(n1322), .B1(LLL3[9]), .Y(n343)
         );
  INVX1 U752 ( .A(n344), .Y(n1012) );
  AOI22X1 U753 ( .A0(n1335), .A1(LLL3[9]), .B0(n1322), .B1(LLL2[9]), .Y(n344)
         );
  INVX1 U754 ( .A(n350), .Y(n1018) );
  AOI22X1 U755 ( .A0(n1333), .A1(LLL7[8]), .B0(n1322), .B1(LLL6[8]), .Y(n350)
         );
  INVX1 U756 ( .A(n351), .Y(n1019) );
  AOI22X1 U757 ( .A0(n1363), .A1(LLL6[8]), .B0(n1322), .B1(LLL5[8]), .Y(n351)
         );
  INVX1 U758 ( .A(n352), .Y(n1020) );
  AOI22X1 U759 ( .A0(n1404), .A1(LLL5[8]), .B0(n1322), .B1(LLL4[8]), .Y(n352)
         );
  INVX1 U760 ( .A(n353), .Y(n1021) );
  AOI22X1 U761 ( .A0(n1330), .A1(LLL4[8]), .B0(n1322), .B1(LLL3[8]), .Y(n353)
         );
  INVX1 U762 ( .A(n354), .Y(n1022) );
  AOI22X1 U763 ( .A0(n1375), .A1(LLL3[8]), .B0(n1322), .B1(LLL2[8]), .Y(n354)
         );
  INVX1 U764 ( .A(n360), .Y(n1028) );
  AOI22X1 U765 ( .A0(n1388), .A1(LLL7[7]), .B0(n1323), .B1(LLL6[7]), .Y(n360)
         );
  INVX1 U766 ( .A(n361), .Y(n1029) );
  AOI22X1 U767 ( .A0(n1371), .A1(LLL6[7]), .B0(n1323), .B1(LLL5[7]), .Y(n361)
         );
  INVX1 U768 ( .A(n362), .Y(n1030) );
  AOI22X1 U769 ( .A0(n1383), .A1(LLL5[7]), .B0(n1323), .B1(LLL4[7]), .Y(n362)
         );
  INVX1 U770 ( .A(n363), .Y(n1031) );
  AOI22X1 U771 ( .A0(n1387), .A1(LLL4[7]), .B0(n1323), .B1(LLL3[7]), .Y(n363)
         );
  INVX1 U772 ( .A(n364), .Y(n1032) );
  AOI22X1 U773 ( .A0(n1330), .A1(LLL3[7]), .B0(n1323), .B1(LLL2[7]), .Y(n364)
         );
  INVX1 U774 ( .A(n370), .Y(n1038) );
  AOI22X1 U775 ( .A0(n1386), .A1(LLL7[6]), .B0(n1323), .B1(LLL6[6]), .Y(n370)
         );
  INVX1 U776 ( .A(n371), .Y(n1039) );
  AOI22X1 U777 ( .A0(n1387), .A1(LLL6[6]), .B0(n1323), .B1(LLL5[6]), .Y(n371)
         );
  INVX1 U778 ( .A(n372), .Y(n1040) );
  AOI22X1 U779 ( .A0(n1336), .A1(LLL5[6]), .B0(n1323), .B1(LLL4[6]), .Y(n372)
         );
  INVX1 U780 ( .A(n373), .Y(n1041) );
  AOI22X1 U781 ( .A0(n1372), .A1(LLL4[6]), .B0(n1323), .B1(LLL3[6]), .Y(n373)
         );
  INVX1 U782 ( .A(n374), .Y(n1042) );
  AOI22X1 U783 ( .A0(n1384), .A1(LLL3[6]), .B0(n1324), .B1(LLL2[6]), .Y(n374)
         );
  INVX1 U784 ( .A(n375), .Y(n1043) );
  AOI22X1 U785 ( .A0(n1376), .A1(LLL2[6]), .B0(n1324), .B1(LLL1[6]), .Y(n375)
         );
  INVX1 U786 ( .A(n380), .Y(n1048) );
  AOI22X1 U787 ( .A0(n1380), .A1(LLL7[5]), .B0(n1324), .B1(LLL6[5]), .Y(n380)
         );
  INVX1 U788 ( .A(n381), .Y(n1049) );
  AOI22X1 U789 ( .A0(n1373), .A1(LLL6[5]), .B0(n1324), .B1(LLL5[5]), .Y(n381)
         );
  INVX1 U790 ( .A(n382), .Y(n1050) );
  AOI22X1 U791 ( .A0(n1381), .A1(LLL5[5]), .B0(n1324), .B1(LLL4[5]), .Y(n382)
         );
  INVX1 U792 ( .A(n383), .Y(n1051) );
  AOI22X1 U793 ( .A0(n1379), .A1(LLL4[5]), .B0(n1324), .B1(LLL3[5]), .Y(n383)
         );
  INVX1 U794 ( .A(n384), .Y(n1052) );
  AOI22X1 U795 ( .A0(n1334), .A1(LLL3[5]), .B0(n1324), .B1(LLL2[5]), .Y(n384)
         );
  INVX1 U796 ( .A(n390), .Y(n1058) );
  AOI22X1 U797 ( .A0(n1330), .A1(LLL7[4]), .B0(n1324), .B1(LLL6[4]), .Y(n390)
         );
  INVX1 U798 ( .A(n391), .Y(n1059) );
  AOI22X1 U799 ( .A0(n1404), .A1(LLL6[4]), .B0(n1324), .B1(LLL5[4]), .Y(n391)
         );
  INVX1 U800 ( .A(n392), .Y(n1060) );
  AOI22X1 U801 ( .A0(n1331), .A1(LLL5[4]), .B0(n1325), .B1(LLL4[4]), .Y(n392)
         );
  INVX1 U802 ( .A(n393), .Y(n1061) );
  AOI22X1 U803 ( .A0(n1332), .A1(LLL4[4]), .B0(n1325), .B1(LLL3[4]), .Y(n393)
         );
  INVX1 U804 ( .A(n394), .Y(n1062) );
  AOI22X1 U805 ( .A0(n1335), .A1(LLL3[4]), .B0(n1325), .B1(LLL2[4]), .Y(n394)
         );
  INVX1 U806 ( .A(n400), .Y(n1068) );
  AOI22X1 U807 ( .A0(n1377), .A1(LLL7[3]), .B0(n1325), .B1(LLL6[3]), .Y(n400)
         );
  INVX1 U808 ( .A(n401), .Y(n1069) );
  AOI22X1 U809 ( .A0(n1360), .A1(LLL6[3]), .B0(n1325), .B1(LLL5[3]), .Y(n401)
         );
  INVX1 U810 ( .A(n402), .Y(n1070) );
  AOI22X1 U811 ( .A0(n1386), .A1(LLL5[3]), .B0(n1325), .B1(LLL4[3]), .Y(n402)
         );
  INVX1 U812 ( .A(n403), .Y(n1071) );
  AOI22X1 U813 ( .A0(n1374), .A1(LLL4[3]), .B0(n1325), .B1(LLL3[3]), .Y(n403)
         );
  INVX1 U814 ( .A(n404), .Y(n1072) );
  AOI22X1 U815 ( .A0(n1351), .A1(LLL3[3]), .B0(n1325), .B1(LLL2[3]), .Y(n404)
         );
  INVX1 U816 ( .A(n410), .Y(n1078) );
  AOI22X1 U817 ( .A0(n1354), .A1(LLL7[2]), .B0(n1326), .B1(LLL6[2]), .Y(n410)
         );
  INVX1 U818 ( .A(n411), .Y(n1079) );
  AOI22X1 U819 ( .A0(n1408), .A1(LLL6[2]), .B0(n1320), .B1(LLL5[2]), .Y(n411)
         );
  INVX1 U820 ( .A(n412), .Y(n1080) );
  AOI22X1 U821 ( .A0(n1342), .A1(LLL5[2]), .B0(n1326), .B1(LLL4[2]), .Y(n412)
         );
  INVX1 U822 ( .A(n413), .Y(n1081) );
  AOI22X1 U823 ( .A0(n1385), .A1(LLL4[2]), .B0(n1326), .B1(LLL3[2]), .Y(n413)
         );
  INVX1 U824 ( .A(n414), .Y(n1082) );
  AOI22X1 U825 ( .A0(n1330), .A1(LLL3[2]), .B0(n1326), .B1(LLL2[2]), .Y(n414)
         );
  INVX1 U826 ( .A(n415), .Y(n1083) );
  AOI22X1 U827 ( .A0(n1365), .A1(LLL2[2]), .B0(n1326), .B1(LLL1[2]), .Y(n415)
         );
  INVX1 U828 ( .A(n420), .Y(n1088) );
  AOI22X1 U829 ( .A0(n1353), .A1(LLL7[1]), .B0(n1327), .B1(LLL6[1]), .Y(n420)
         );
  INVX1 U830 ( .A(n421), .Y(n1089) );
  AOI22X1 U831 ( .A0(n1359), .A1(LLL6[1]), .B0(n1326), .B1(LLL5[1]), .Y(n421)
         );
  INVX1 U832 ( .A(n422), .Y(n1090) );
  AOI22X1 U833 ( .A0(n1346), .A1(LLL5[1]), .B0(n1327), .B1(LLL4[1]), .Y(n422)
         );
  INVX1 U834 ( .A(n423), .Y(n1091) );
  AOI22X1 U835 ( .A0(n1362), .A1(LLL4[1]), .B0(n1327), .B1(LLL3[1]), .Y(n423)
         );
  INVX1 U836 ( .A(n424), .Y(n1092) );
  AOI22X1 U837 ( .A0(n1364), .A1(LLL3[1]), .B0(n1328), .B1(LLL2[1]), .Y(n424)
         );
  INVX1 U838 ( .A(n425), .Y(n1093) );
  AOI22X1 U839 ( .A0(n1366), .A1(LLL2[1]), .B0(n1327), .B1(LLL1[1]), .Y(n425)
         );
  INVX1 U840 ( .A(n430), .Y(n1098) );
  AOI22X1 U841 ( .A0(n1331), .A1(LLL7[0]), .B0(n1328), .B1(LLL6[0]), .Y(n430)
         );
  INVX1 U842 ( .A(n431), .Y(n1099) );
  AOI22X1 U843 ( .A0(n1405), .A1(LLL6[0]), .B0(n1326), .B1(LLL5[0]), .Y(n431)
         );
  INVX1 U844 ( .A(n432), .Y(n1100) );
  AOI22X1 U845 ( .A0(n1347), .A1(LLL5[0]), .B0(n1328), .B1(LLL4[0]), .Y(n432)
         );
  INVX1 U846 ( .A(n433), .Y(n1101) );
  AOI22X1 U847 ( .A0(n1365), .A1(LLL4[0]), .B0(n1326), .B1(LLL3[0]), .Y(n433)
         );
  INVX1 U848 ( .A(n434), .Y(n1102) );
  AOI22X1 U849 ( .A0(n1345), .A1(LLL3[0]), .B0(n644), .B1(LLL2[0]), .Y(n434)
         );
  INVX1 U850 ( .A(n435), .Y(n1103) );
  AOI22X1 U851 ( .A0(n1367), .A1(LLL2[0]), .B0(n1327), .B1(LLL1[0]), .Y(n435)
         );
  INVX1 U852 ( .A(n438), .Y(n1106) );
  AOI22X1 U853 ( .A0(n650), .A1(U6[12]), .B0(n1369), .B1(U7[12]), .Y(n438) );
  INVX1 U854 ( .A(n439), .Y(n1107) );
  AOI22X1 U855 ( .A0(n652), .A1(U5[12]), .B0(n1369), .B1(U6[12]), .Y(n439) );
  INVX1 U856 ( .A(n440), .Y(n1108) );
  AOI22X1 U857 ( .A0(n649), .A1(U4[12]), .B0(n1368), .B1(U5[12]), .Y(n440) );
  INVX1 U858 ( .A(n441), .Y(n1109) );
  AOI22X1 U859 ( .A0(n649), .A1(U3[12]), .B0(n1364), .B1(U4[12]), .Y(n441) );
  INVX1 U860 ( .A(n442), .Y(n1110) );
  AOI22X1 U861 ( .A0(n649), .A1(U2[12]), .B0(n1380), .B1(U3[12]), .Y(n442) );
  INVX1 U862 ( .A(n443), .Y(n1111) );
  AOI22X1 U863 ( .A0(n649), .A1(U1[12]), .B0(n1374), .B1(U2[12]), .Y(n443) );
  INVX1 U864 ( .A(n444), .Y(n1112) );
  AOI22X1 U865 ( .A0(n649), .A1(Uout[12]), .B0(n1384), .B1(U1[12]), .Y(n444)
         );
  INVX1 U866 ( .A(n447), .Y(n1115) );
  AOI22X1 U867 ( .A0(n649), .A1(U6[11]), .B0(n1408), .B1(U7[11]), .Y(n447) );
  INVX1 U868 ( .A(n448), .Y(n1116) );
  AOI22X1 U869 ( .A0(n649), .A1(U5[11]), .B0(n1349), .B1(U6[11]), .Y(n448) );
  INVX1 U870 ( .A(n449), .Y(n1117) );
  AOI22X1 U871 ( .A0(n656), .A1(U4[11]), .B0(n1367), .B1(U5[11]), .Y(n449) );
  INVX1 U872 ( .A(n450), .Y(n1118) );
  AOI22X1 U873 ( .A0(n806), .A1(U3[11]), .B0(n1358), .B1(U4[11]), .Y(n450) );
  INVX1 U874 ( .A(n451), .Y(n1119) );
  AOI22X1 U875 ( .A0(n806), .A1(U2[11]), .B0(n1360), .B1(U3[11]), .Y(n451) );
  INVX1 U876 ( .A(n452), .Y(n1120) );
  AOI22X1 U877 ( .A0(n806), .A1(U1[11]), .B0(n1346), .B1(U2[11]), .Y(n452) );
  INVX1 U878 ( .A(n453), .Y(n1121) );
  AOI22X1 U879 ( .A0(n806), .A1(Uout[11]), .B0(n1366), .B1(U1[11]), .Y(n453)
         );
  INVX1 U880 ( .A(n456), .Y(n1124) );
  AOI22X1 U881 ( .A0(n798), .A1(U6[10]), .B0(n1338), .B1(U7[10]), .Y(n456) );
  INVX1 U882 ( .A(n457), .Y(n1125) );
  AOI22X1 U883 ( .A0(n798), .A1(U5[10]), .B0(n1374), .B1(U6[10]), .Y(n457) );
  INVX1 U884 ( .A(n458), .Y(n1126) );
  AOI22X1 U885 ( .A0(n798), .A1(U4[10]), .B0(n1359), .B1(U5[10]), .Y(n458) );
  INVX1 U886 ( .A(n459), .Y(n1127) );
  AOI22X1 U887 ( .A0(n798), .A1(U3[10]), .B0(n1350), .B1(U4[10]), .Y(n459) );
  INVX1 U888 ( .A(n460), .Y(n1128) );
  AOI22X1 U889 ( .A0(n798), .A1(U2[10]), .B0(n1355), .B1(U3[10]), .Y(n460) );
  INVX1 U890 ( .A(n461), .Y(n1129) );
  AOI22X1 U891 ( .A0(n798), .A1(U1[10]), .B0(n1367), .B1(U2[10]), .Y(n461) );
  INVX1 U892 ( .A(n462), .Y(n1130) );
  AOI22X1 U893 ( .A0(n798), .A1(Uout[10]), .B0(n1363), .B1(U1[10]), .Y(n462)
         );
  INVX1 U894 ( .A(n465), .Y(n1133) );
  AOI22X1 U895 ( .A0(n790), .A1(U6[9]), .B0(n1401), .B1(U7[9]), .Y(n465) );
  INVX1 U896 ( .A(n466), .Y(n1134) );
  AOI22X1 U897 ( .A0(n790), .A1(U5[9]), .B0(n1352), .B1(U6[9]), .Y(n466) );
  INVX1 U898 ( .A(n467), .Y(n1135) );
  AOI22X1 U899 ( .A0(n790), .A1(U4[9]), .B0(n1380), .B1(U5[9]), .Y(n467) );
  INVX1 U900 ( .A(n468), .Y(n1136) );
  AOI22X1 U901 ( .A0(n790), .A1(U3[9]), .B0(n1368), .B1(U4[9]), .Y(n468) );
  INVX1 U902 ( .A(n469), .Y(n1137) );
  AOI22X1 U903 ( .A0(n790), .A1(U2[9]), .B0(n1362), .B1(U3[9]), .Y(n469) );
  INVX1 U904 ( .A(n470), .Y(n1138) );
  AOI22X1 U905 ( .A0(n790), .A1(U1[9]), .B0(n1359), .B1(U2[9]), .Y(n470) );
  INVX1 U906 ( .A(n471), .Y(n1139) );
  AOI22X1 U907 ( .A0(n790), .A1(Uout[9]), .B0(n1350), .B1(U1[9]), .Y(n471) );
  INVX1 U908 ( .A(n474), .Y(n1142) );
  AOI22X1 U909 ( .A0(n790), .A1(U6[8]), .B0(n1353), .B1(U7[8]), .Y(n474) );
  INVX1 U910 ( .A(n475), .Y(n1143) );
  AOI22X1 U911 ( .A0(n782), .A1(U5[8]), .B0(n1387), .B1(U6[8]), .Y(n475) );
  INVX1 U912 ( .A(n476), .Y(n1144) );
  AOI22X1 U913 ( .A0(n782), .A1(U4[8]), .B0(n1370), .B1(U5[8]), .Y(n476) );
  INVX1 U914 ( .A(n477), .Y(n1145) );
  AOI22X1 U915 ( .A0(n782), .A1(U3[8]), .B0(n1401), .B1(U4[8]), .Y(n477) );
  INVX1 U916 ( .A(n478), .Y(n1146) );
  AOI22X1 U917 ( .A0(n782), .A1(U2[8]), .B0(n1361), .B1(U3[8]), .Y(n478) );
  INVX1 U918 ( .A(n479), .Y(n1147) );
  AOI22X1 U919 ( .A0(n782), .A1(U1[8]), .B0(n1354), .B1(U2[8]), .Y(n479) );
  INVX1 U920 ( .A(n480), .Y(n1148) );
  AOI22X1 U921 ( .A0(n782), .A1(Uout[8]), .B0(n1382), .B1(U1[8]), .Y(n480) );
  INVX1 U922 ( .A(n483), .Y(n1151) );
  AOI22X1 U923 ( .A0(n782), .A1(U6[7]), .B0(n1383), .B1(U7[7]), .Y(n483) );
  INVX1 U924 ( .A(n484), .Y(n1152) );
  AOI22X1 U925 ( .A0(n782), .A1(U5[7]), .B0(n1380), .B1(U6[7]), .Y(n484) );
  INVX1 U926 ( .A(n485), .Y(n1153) );
  AOI22X1 U927 ( .A0(n670), .A1(U4[7]), .B0(n1337), .B1(U5[7]), .Y(n485) );
  INVX1 U928 ( .A(n486), .Y(n1154) );
  AOI22X1 U929 ( .A0(n670), .A1(U3[7]), .B0(n1366), .B1(U4[7]), .Y(n486) );
  INVX1 U930 ( .A(n487), .Y(n1155) );
  AOI22X1 U931 ( .A0(n670), .A1(U2[7]), .B0(n1381), .B1(U3[7]), .Y(n487) );
  INVX1 U932 ( .A(n488), .Y(n1156) );
  AOI22X1 U933 ( .A0(n1004), .A1(U1[7]), .B0(n1348), .B1(U2[7]), .Y(n488) );
  INVX1 U934 ( .A(n489), .Y(n1157) );
  AOI22X1 U935 ( .A0(n670), .A1(Uout[7]), .B0(n1344), .B1(U1[7]), .Y(n489) );
  INVX1 U936 ( .A(n492), .Y(n1160) );
  AOI22X1 U937 ( .A0(n670), .A1(U6[6]), .B0(n1405), .B1(U7[6]), .Y(n492) );
  INVX1 U938 ( .A(n493), .Y(n1161) );
  AOI22X1 U939 ( .A0(n670), .A1(U5[6]), .B0(n1378), .B1(U6[6]), .Y(n493) );
  INVX1 U940 ( .A(n494), .Y(n1162) );
  AOI22X1 U941 ( .A0(n670), .A1(U4[6]), .B0(n1381), .B1(U5[6]), .Y(n494) );
  INVX1 U942 ( .A(n495), .Y(n1163) );
  AOI22X1 U943 ( .A0(n670), .A1(U3[6]), .B0(n1349), .B1(U4[6]), .Y(n495) );
  INVX1 U944 ( .A(n496), .Y(n1164) );
  AOI22X1 U945 ( .A0(n669), .A1(U2[6]), .B0(n1377), .B1(U3[6]), .Y(n496) );
  INVX1 U946 ( .A(n497), .Y(n1165) );
  AOI22X1 U947 ( .A0(n669), .A1(U1[6]), .B0(n1386), .B1(U2[6]), .Y(n497) );
  INVX1 U948 ( .A(n498), .Y(n1166) );
  AOI22X1 U949 ( .A0(n669), .A1(Uout[6]), .B0(n1341), .B1(U1[6]), .Y(n498) );
  INVX1 U950 ( .A(n501), .Y(n1169) );
  AOI22X1 U951 ( .A0(n669), .A1(U6[5]), .B0(n1350), .B1(U7[5]), .Y(n501) );
  INVX1 U952 ( .A(n502), .Y(n1170) );
  AOI22X1 U953 ( .A0(n669), .A1(U5[5]), .B0(n1380), .B1(U6[5]), .Y(n502) );
  INVX1 U954 ( .A(n503), .Y(n1171) );
  AOI22X1 U955 ( .A0(n669), .A1(U4[5]), .B0(n1345), .B1(U5[5]), .Y(n503) );
  INVX1 U956 ( .A(n504), .Y(n1172) );
  AOI22X1 U957 ( .A0(n669), .A1(U3[5]), .B0(n1342), .B1(U4[5]), .Y(n504) );
  INVX1 U958 ( .A(n505), .Y(n1173) );
  AOI22X1 U959 ( .A0(n669), .A1(U2[5]), .B0(n1343), .B1(U3[5]), .Y(n505) );
  INVX1 U960 ( .A(n506), .Y(n1174) );
  AOI22X1 U961 ( .A0(n668), .A1(U1[5]), .B0(n1347), .B1(U2[5]), .Y(n506) );
  INVX1 U962 ( .A(n507), .Y(n1175) );
  AOI22X1 U963 ( .A0(n668), .A1(Uout[5]), .B0(n1368), .B1(U1[5]), .Y(n507) );
  INVX1 U964 ( .A(n510), .Y(n1178) );
  AOI22X1 U965 ( .A0(n668), .A1(U6[4]), .B0(n1338), .B1(U7[4]), .Y(n510) );
  INVX1 U966 ( .A(n511), .Y(n1179) );
  AOI22X1 U967 ( .A0(n668), .A1(U5[4]), .B0(n1367), .B1(U6[4]), .Y(n511) );
  INVX1 U968 ( .A(n512), .Y(n1180) );
  AOI22X1 U969 ( .A0(n668), .A1(U4[4]), .B0(n1359), .B1(U5[4]), .Y(n512) );
  INVX1 U970 ( .A(n513), .Y(n1181) );
  AOI22X1 U971 ( .A0(n668), .A1(U3[4]), .B0(n1352), .B1(U4[4]), .Y(n513) );
  INVX1 U972 ( .A(n514), .Y(n1182) );
  AOI22X1 U973 ( .A0(n668), .A1(U2[4]), .B0(n1365), .B1(U3[4]), .Y(n514) );
  INVX1 U974 ( .A(n515), .Y(n1183) );
  AOI22X1 U975 ( .A0(n667), .A1(U1[4]), .B0(n1353), .B1(U2[4]), .Y(n515) );
  INVX1 U976 ( .A(n516), .Y(n1184) );
  AOI22X1 U977 ( .A0(n667), .A1(Uout[4]), .B0(n1357), .B1(U1[4]), .Y(n516) );
  INVX1 U978 ( .A(n519), .Y(n1187) );
  AOI22X1 U979 ( .A0(n667), .A1(U6[3]), .B0(n1351), .B1(U7[3]), .Y(n519) );
  INVX1 U980 ( .A(n520), .Y(n1188) );
  AOI22X1 U981 ( .A0(n667), .A1(U5[3]), .B0(n1346), .B1(U6[3]), .Y(n520) );
  INVX1 U982 ( .A(n521), .Y(n1189) );
  AOI22X1 U983 ( .A0(n667), .A1(U4[3]), .B0(n1355), .B1(U5[3]), .Y(n521) );
  INVX1 U984 ( .A(n522), .Y(n1190) );
  AOI22X1 U985 ( .A0(n667), .A1(U3[3]), .B0(n1369), .B1(U4[3]), .Y(n522) );
  INVX1 U986 ( .A(n523), .Y(n1191) );
  AOI22X1 U987 ( .A0(n667), .A1(U2[3]), .B0(n1340), .B1(U3[3]), .Y(n523) );
  INVX1 U988 ( .A(n524), .Y(n1192) );
  AOI22X1 U989 ( .A0(n667), .A1(U1[3]), .B0(n1408), .B1(U2[3]), .Y(n524) );
  INVX1 U990 ( .A(n528), .Y(n1196) );
  AOI22X1 U991 ( .A0(n666), .A1(U6[2]), .B0(n1349), .B1(U7[2]), .Y(n528) );
  INVX1 U992 ( .A(n529), .Y(n1197) );
  AOI22X1 U993 ( .A0(n666), .A1(U5[2]), .B0(n1348), .B1(U6[2]), .Y(n529) );
  INVX1 U994 ( .A(n530), .Y(n1198) );
  AOI22X1 U995 ( .A0(n666), .A1(U4[2]), .B0(n1344), .B1(U5[2]), .Y(n530) );
  INVX1 U996 ( .A(n531), .Y(n1199) );
  AOI22X1 U997 ( .A0(n666), .A1(U3[2]), .B0(n1362), .B1(U4[2]), .Y(n531) );
  INVX1 U998 ( .A(n532), .Y(n1200) );
  AOI22X1 U999 ( .A0(n666), .A1(U2[2]), .B0(n1356), .B1(U3[2]), .Y(n532) );
  INVX1 U1000 ( .A(n533), .Y(n1201) );
  AOI22X1 U1001 ( .A0(n666), .A1(U1[2]), .B0(n1382), .B1(U2[2]), .Y(n533) );
  INVX1 U1002 ( .A(n537), .Y(n1205) );
  AOI22X1 U1003 ( .A0(n665), .A1(U6[1]), .B0(n1364), .B1(U7[1]), .Y(n537) );
  INVX1 U1004 ( .A(n538), .Y(n1206) );
  AOI22X1 U1005 ( .A0(n665), .A1(U5[1]), .B0(n1365), .B1(U6[1]), .Y(n538) );
  INVX1 U1006 ( .A(n539), .Y(n1207) );
  AOI22X1 U1007 ( .A0(n665), .A1(U4[1]), .B0(n1400), .B1(U5[1]), .Y(n539) );
  INVX1 U1008 ( .A(n540), .Y(n1208) );
  AOI22X1 U1009 ( .A0(n665), .A1(U3[1]), .B0(n1357), .B1(U4[1]), .Y(n540) );
  INVX1 U1010 ( .A(n541), .Y(n1209) );
  AOI22X1 U1011 ( .A0(n665), .A1(U2[1]), .B0(n1360), .B1(U3[1]), .Y(n541) );
  INVX1 U1012 ( .A(n542), .Y(n1210) );
  AOI22X1 U1013 ( .A0(n665), .A1(U1[1]), .B0(n1408), .B1(U2[1]), .Y(n542) );
  INVX1 U1014 ( .A(n543), .Y(n1211) );
  AOI22X1 U1015 ( .A0(n665), .A1(Uout[1]), .B0(n1366), .B1(U1[1]), .Y(n543) );
  INVX1 U1016 ( .A(n546), .Y(n1214) );
  AOI22X1 U1017 ( .A0(n664), .A1(U6[0]), .B0(n1370), .B1(U7[0]), .Y(n546) );
  INVX1 U1018 ( .A(n547), .Y(n1215) );
  AOI22X1 U1019 ( .A0(n664), .A1(U5[0]), .B0(n1402), .B1(U6[0]), .Y(n547) );
  INVX1 U1020 ( .A(n548), .Y(n1216) );
  AOI22X1 U1021 ( .A0(n664), .A1(U4[0]), .B0(n1385), .B1(U5[0]), .Y(n548) );
  INVX1 U1022 ( .A(n549), .Y(n1217) );
  AOI22X1 U1023 ( .A0(n664), .A1(U3[0]), .B0(n1367), .B1(U4[0]), .Y(n549) );
  INVX1 U1024 ( .A(n550), .Y(n1218) );
  AOI22X1 U1025 ( .A0(n664), .A1(U2[0]), .B0(n1390), .B1(U3[0]), .Y(n550) );
  INVX1 U1026 ( .A(n551), .Y(n1219) );
  AOI22X1 U1027 ( .A0(n664), .A1(U1[0]), .B0(n1340), .B1(U2[0]), .Y(n551) );
  INVX1 U1028 ( .A(n552), .Y(n1220) );
  AOI22X1 U1029 ( .A0(n664), .A1(Uout[0]), .B0(n1377), .B1(U1[0]), .Y(n552) );
  INVX1 U1030 ( .A(n14), .Y(n681) );
  AOI22X1 U1031 ( .A0(n1333), .A1(DR1[4]), .B0(deg_Ro[4]), .B1(n1054), .Y(n14)
         );
  INVX1 U1032 ( .A(n22), .Y(n689) );
  AOI22X1 U1033 ( .A0(n1340), .A1(DR1[3]), .B0(deg_Ro[3]), .B1(n1054), .Y(n22)
         );
  INVX1 U1034 ( .A(n30), .Y(n697) );
  AOI22X1 U1035 ( .A0(n1333), .A1(DR1[2]), .B0(deg_Ro[2]), .B1(n1034), .Y(n30)
         );
  INVX1 U1036 ( .A(n38), .Y(n705) );
  AOI22X1 U1037 ( .A0(n1331), .A1(DR1[1]), .B0(deg_Ro[1]), .B1(n1054), .Y(n38)
         );
  INVX1 U1038 ( .A(n46), .Y(n713) );
  AOI22X1 U1039 ( .A0(n1333), .A1(DR1[0]), .B0(deg_Ro[0]), .B1(n1046), .Y(n46)
         );
  INVX1 U1040 ( .A(n54), .Y(n721) );
  AOI22X1 U1041 ( .A0(n1381), .A1(DQ1[4]), .B0(deg_Qo[4]), .B1(n1054), .Y(n54)
         );
  INVX1 U1042 ( .A(n62), .Y(n729) );
  AOI22X1 U1043 ( .A0(n1383), .A1(DQ1[3]), .B0(deg_Qo[3]), .B1(n1034), .Y(n62)
         );
  INVX1 U1044 ( .A(n70), .Y(n737) );
  AOI22X1 U1045 ( .A0(n1336), .A1(DQ1[2]), .B0(deg_Qo[2]), .B1(n1046), .Y(n70)
         );
  INVX1 U1046 ( .A(n78), .Y(n745) );
  AOI22X1 U1047 ( .A0(n1387), .A1(DQ1[1]), .B0(deg_Qo[1]), .B1(n1034), .Y(n78)
         );
  INVX1 U1048 ( .A(n86), .Y(n753) );
  AOI22X1 U1049 ( .A0(n1390), .A1(DQ1[0]), .B0(deg_Qo[0]), .B1(n1046), .Y(n86)
         );
  INVX1 U1050 ( .A(n210), .Y(n878) );
  AOI22X1 U1051 ( .A0(n1356), .A1(Q1[12]), .B0(Qout[12]), .B1(n1046), .Y(n210)
         );
  INVX1 U1052 ( .A(n218), .Y(n886) );
  AOI22X1 U1053 ( .A0(n1347), .A1(Q1[11]), .B0(Qout[11]), .B1(n1034), .Y(n218)
         );
  INVX1 U1054 ( .A(n226), .Y(n894) );
  AOI22X1 U1055 ( .A0(n1355), .A1(Q1[10]), .B0(Qout[10]), .B1(n1046), .Y(n226)
         );
  INVX1 U1056 ( .A(n234), .Y(n902) );
  AOI22X1 U1057 ( .A0(n1331), .A1(Q1[9]), .B0(Qout[9]), .B1(n1054), .Y(n234)
         );
  INVX1 U1058 ( .A(n242), .Y(n910) );
  AOI22X1 U1059 ( .A0(n1353), .A1(Q1[8]), .B0(Qout[8]), .B1(n1046), .Y(n242)
         );
  INVX1 U1060 ( .A(n250), .Y(n918) );
  AOI22X1 U1061 ( .A0(n1376), .A1(Q1[7]), .B0(Qout[7]), .B1(n1046), .Y(n250)
         );
  INVX1 U1062 ( .A(n258), .Y(n926) );
  AOI22X1 U1063 ( .A0(n1331), .A1(Q1[6]), .B0(Qout[6]), .B1(n1054), .Y(n258)
         );
  INVX1 U1064 ( .A(n266), .Y(n934) );
  AOI22X1 U1065 ( .A0(n1370), .A1(Q1[5]), .B0(Qout[5]), .B1(n1056), .Y(n266)
         );
  INVX1 U1066 ( .A(n274), .Y(n942) );
  AOI22X1 U1067 ( .A0(n1348), .A1(Q1[4]), .B0(Qout[4]), .B1(n1054), .Y(n274)
         );
  INVX1 U1068 ( .A(n282), .Y(n950) );
  AOI22X1 U1069 ( .A0(n1363), .A1(Q1[3]), .B0(Qout[3]), .B1(n1054), .Y(n282)
         );
  INVX1 U1070 ( .A(n290), .Y(n958) );
  AOI22X1 U1071 ( .A0(n1352), .A1(Q1[2]), .B0(Qout[2]), .B1(n1056), .Y(n290)
         );
  INVX1 U1072 ( .A(n298), .Y(n966) );
  AOI22X1 U1073 ( .A0(n1367), .A1(Q1[1]), .B0(Qout[1]), .B1(n1066), .Y(n298)
         );
  INVX1 U1074 ( .A(n306), .Y(n974) );
  AOI22X1 U1075 ( .A0(n1350), .A1(Q1[0]), .B0(Qout[0]), .B1(n1314), .Y(n306)
         );
  INVX1 U1076 ( .A(n325), .Y(n993) );
  AOI22X1 U1077 ( .A0(n1332), .A1(LLL2[11]), .B0(n1320), .B1(LLL1[11]), .Y(
        n325) );
  INVX1 U1078 ( .A(n335), .Y(n1003) );
  AOI22X1 U1079 ( .A0(n1330), .A1(LLL2[10]), .B0(n1321), .B1(LLL1[10]), .Y(
        n335) );
  INVX1 U1080 ( .A(n345), .Y(n1013) );
  AOI22X1 U1081 ( .A0(n1334), .A1(LLL2[9]), .B0(n1322), .B1(LLL1[9]), .Y(n345)
         );
  INVX1 U1082 ( .A(n355), .Y(n1023) );
  AOI22X1 U1083 ( .A0(n1379), .A1(LLL2[8]), .B0(n1322), .B1(LLL1[8]), .Y(n355)
         );
  INVX1 U1084 ( .A(n365), .Y(n1033) );
  AOI22X1 U1085 ( .A0(n1333), .A1(LLL2[7]), .B0(n1323), .B1(LLL1[7]), .Y(n365)
         );
  INVX1 U1086 ( .A(n385), .Y(n1053) );
  AOI22X1 U1087 ( .A0(n1332), .A1(LLL2[5]), .B0(n1324), .B1(LLL1[5]), .Y(n385)
         );
  INVX1 U1088 ( .A(n571), .Y(n1240) );
  AOI22X1 U1089 ( .A0(n1374), .A1(count[9]), .B0(N185), .B1(n1064), .Y(n571)
         );
  INVX1 U1090 ( .A(n576), .Y(n1245) );
  AOI22X1 U1091 ( .A0(n1337), .A1(count[4]), .B0(N180), .B1(n1056), .Y(n576)
         );
  INVX1 U1092 ( .A(n578), .Y(n1247) );
  AOI22X1 U1093 ( .A0(n1340), .A1(count[2]), .B0(N178), .B1(n1064), .Y(n578)
         );
  INVX1 U1094 ( .A(n580), .Y(n1249) );
  AOI22X1 U1095 ( .A0(n1340), .A1(count[0]), .B0(N176), .B1(n1056), .Y(n580)
         );
  INVX1 U1096 ( .A(n581), .Y(n1250) );
  AOI22X1 U1097 ( .A0(Uin_reg[0]), .A1(n1363), .B0(Uin[0]), .B1(n1066), .Y(
        n581) );
  INVX1 U1098 ( .A(n582), .Y(n1251) );
  AOI22X1 U1099 ( .A0(Uin_reg[1]), .A1(n1339), .B0(Uin[1]), .B1(n1066), .Y(
        n582) );
  INVX1 U1100 ( .A(n583), .Y(n1252) );
  AOI22X1 U1101 ( .A0(Uin_reg[2]), .A1(n1369), .B0(Uin[2]), .B1(n1064), .Y(
        n583) );
  INVX1 U1102 ( .A(n584), .Y(n1253) );
  AOI22X1 U1103 ( .A0(Uin_reg[3]), .A1(n1386), .B0(Uin[3]), .B1(n1066), .Y(
        n584) );
  INVX1 U1104 ( .A(n585), .Y(n1254) );
  AOI22X1 U1105 ( .A0(Uin_reg[4]), .A1(n1403), .B0(Uin[4]), .B1(n1066), .Y(
        n585) );
  INVX1 U1106 ( .A(n586), .Y(n1255) );
  AOI22X1 U1107 ( .A0(Uin_reg[5]), .A1(n1403), .B0(Uin[5]), .B1(n1066), .Y(
        n586) );
  INVX1 U1108 ( .A(n587), .Y(n1256) );
  AOI22X1 U1109 ( .A0(Uin_reg[6]), .A1(n1358), .B0(Uin[6]), .B1(n1064), .Y(
        n587) );
  INVX1 U1110 ( .A(n588), .Y(n1257) );
  AOI22X1 U1111 ( .A0(Uin_reg[7]), .A1(n1344), .B0(Uin[7]), .B1(n1064), .Y(
        n588) );
  INVX1 U1112 ( .A(n589), .Y(n1258) );
  AOI22X1 U1113 ( .A0(Uin_reg[8]), .A1(n1333), .B0(Uin[8]), .B1(n1074), .Y(
        n589) );
  INVX1 U1114 ( .A(n590), .Y(n1259) );
  AOI22X1 U1115 ( .A0(Uin_reg[9]), .A1(n1405), .B0(Uin[9]), .B1(n1074), .Y(
        n590) );
  INVX1 U1116 ( .A(n591), .Y(n1260) );
  AOI22X1 U1117 ( .A0(Uin_reg[10]), .A1(n1368), .B0(Uin[10]), .B1(n1066), .Y(
        n591) );
  INVX1 U1118 ( .A(n592), .Y(n1261) );
  AOI22X1 U1119 ( .A0(Uin_reg[11]), .A1(n1388), .B0(Uin[11]), .B1(n1056), .Y(
        n592) );
  INVX1 U1120 ( .A(n593), .Y(n1262) );
  AOI22X1 U1121 ( .A0(Uin_reg[12]), .A1(n1337), .B0(Uin[12]), .B1(n1074), .Y(
        n593) );
  INVX1 U1122 ( .A(n607), .Y(n1276) );
  AOI22X1 U1123 ( .A0(Qin_reg[0]), .A1(n1361), .B0(Qin[0]), .B1(n1066), .Y(
        n607) );
  INVX1 U1124 ( .A(n608), .Y(n1277) );
  AOI22X1 U1125 ( .A0(Qin_reg[1]), .A1(n1384), .B0(Qin[1]), .B1(n1074), .Y(
        n608) );
  INVX1 U1126 ( .A(n609), .Y(n1278) );
  AOI22X1 U1127 ( .A0(Qin_reg[2]), .A1(n1372), .B0(Qin[2]), .B1(n1064), .Y(
        n609) );
  INVX1 U1128 ( .A(n610), .Y(n1279) );
  AOI22X1 U1129 ( .A0(Qin_reg[3]), .A1(n1379), .B0(Qin[3]), .B1(n1074), .Y(
        n610) );
  INVX1 U1130 ( .A(n611), .Y(n1280) );
  AOI22X1 U1131 ( .A0(Qin_reg[4]), .A1(n1405), .B0(Qin[4]), .B1(n1066), .Y(
        n611) );
  INVX1 U1132 ( .A(n612), .Y(n1281) );
  AOI22X1 U1133 ( .A0(Qin_reg[5]), .A1(n1384), .B0(Qin[5]), .B1(n1314), .Y(
        n612) );
  INVX1 U1134 ( .A(n613), .Y(n1282) );
  AOI22X1 U1135 ( .A0(Qin_reg[6]), .A1(n1331), .B0(Qin[6]), .B1(n1314), .Y(
        n613) );
  INVX1 U1136 ( .A(n614), .Y(n1283) );
  AOI22X1 U1137 ( .A0(Qin_reg[7]), .A1(n1355), .B0(Qin[7]), .B1(n1074), .Y(
        n614) );
  INVX1 U1138 ( .A(n615), .Y(n1284) );
  AOI22X1 U1139 ( .A0(Qin_reg[8]), .A1(n1349), .B0(Qin[8]), .B1(n1314), .Y(
        n615) );
  INVX1 U1140 ( .A(n616), .Y(n1285) );
  AOI22X1 U1141 ( .A0(Qin_reg[9]), .A1(n1343), .B0(Qin[9]), .B1(n1314), .Y(
        n616) );
  INVX1 U1142 ( .A(n617), .Y(n1286) );
  AOI22X1 U1143 ( .A0(Qin_reg[10]), .A1(n1348), .B0(Qin[10]), .B1(n1074), .Y(
        n617) );
  INVX1 U1144 ( .A(n618), .Y(n1287) );
  AOI22X1 U1145 ( .A0(Qin_reg[11]), .A1(n1376), .B0(Qin[11]), .B1(n1074), .Y(
        n618) );
  INVX1 U1146 ( .A(n619), .Y(n1288) );
  AOI22X1 U1147 ( .A0(Qin_reg[12]), .A1(n1374), .B0(Qin[12]), .B1(n1314), .Y(
        n619) );
  INVX1 U1148 ( .A(n620), .Y(n1289) );
  AOI22X1 U1149 ( .A0(Rin_reg[0]), .A1(n1342), .B0(Rin[0]), .B1(n1315), .Y(
        n620) );
  INVX1 U1150 ( .A(n621), .Y(n1290) );
  AOI22X1 U1151 ( .A0(Rin_reg[1]), .A1(n1373), .B0(Rin[1]), .B1(n1315), .Y(
        n621) );
  INVX1 U1152 ( .A(n622), .Y(n1291) );
  AOI22X1 U1153 ( .A0(Rin_reg[2]), .A1(n1371), .B0(Rin[2]), .B1(n1314), .Y(
        n622) );
  INVX1 U1154 ( .A(n623), .Y(n1292) );
  AOI22X1 U1155 ( .A0(Rin_reg[3]), .A1(n1337), .B0(Rin[3]), .B1(n1315), .Y(
        n623) );
  INVX1 U1156 ( .A(n624), .Y(n1293) );
  AOI22X1 U1157 ( .A0(Rin_reg[4]), .A1(n1376), .B0(Rin[4]), .B1(n1315), .Y(
        n624) );
  INVX1 U1158 ( .A(n625), .Y(n1294) );
  AOI22X1 U1159 ( .A0(Rin_reg[5]), .A1(n1371), .B0(Rin[5]), .B1(n1315), .Y(
        n625) );
  INVX1 U1160 ( .A(n626), .Y(n1295) );
  AOI22X1 U1161 ( .A0(Rin_reg[6]), .A1(n1354), .B0(Rin[6]), .B1(n1074), .Y(
        n626) );
  INVX1 U1162 ( .A(n627), .Y(n1296) );
  AOI22X1 U1163 ( .A0(Rin_reg[7]), .A1(n1370), .B0(Rin[7]), .B1(n1315), .Y(
        n627) );
  INVX1 U1164 ( .A(n628), .Y(n1297) );
  AOI22X1 U1165 ( .A0(Rin_reg[8]), .A1(n1354), .B0(Rin[8]), .B1(n1314), .Y(
        n628) );
  INVX1 U1166 ( .A(n629), .Y(n1298) );
  AOI22X1 U1167 ( .A0(Rin_reg[9]), .A1(n1343), .B0(Rin[9]), .B1(n1314), .Y(
        n629) );
  INVX1 U1168 ( .A(n630), .Y(n1299) );
  AOI22X1 U1169 ( .A0(Rin_reg[10]), .A1(n1352), .B0(Rin[10]), .B1(n1315), .Y(
        n630) );
  INVX1 U1170 ( .A(n631), .Y(n1300) );
  AOI22X1 U1171 ( .A0(Rin_reg[11]), .A1(n1385), .B0(Rin[11]), .B1(n1316), .Y(
        n631) );
  INVX1 U1172 ( .A(n632), .Y(n1301) );
  AOI22X1 U1173 ( .A0(Rin_reg[12]), .A1(n1347), .B0(Rin[12]), .B1(n1314), .Y(
        n632) );
  INVX1 U1174 ( .A(n633), .Y(n1304) );
  AOI22X1 U1175 ( .A0(dQ_reg[0]), .A1(n1351), .B0(deg_Qi[0]), .B1(n1316), .Y(
        n633) );
  INVX1 U1176 ( .A(n634), .Y(n1305) );
  AOI22X1 U1177 ( .A0(dQ_reg[1]), .A1(n1358), .B0(deg_Qi[1]), .B1(n1315), .Y(
        n634) );
  INVX1 U1178 ( .A(n635), .Y(n1306) );
  AOI22X1 U1179 ( .A0(dQ_reg[2]), .A1(n1357), .B0(deg_Qi[2]), .B1(n1316), .Y(
        n635) );
  INVX1 U1180 ( .A(n636), .Y(n1307) );
  AOI22X1 U1181 ( .A0(dQ_reg[3]), .A1(n1354), .B0(deg_Qi[3]), .B1(n1315), .Y(
        n636) );
  INVX1 U1182 ( .A(n637), .Y(n1308) );
  AOI22X1 U1183 ( .A0(dQ_reg[4]), .A1(n1356), .B0(deg_Qi[4]), .B1(n1316), .Y(
        n637) );
  INVX1 U1184 ( .A(n638), .Y(n1309) );
  AOI22X1 U1185 ( .A0(dR_reg[0]), .A1(n1353), .B0(deg_Ri[0]), .B1(n1316), .Y(
        n638) );
  INVX1 U1186 ( .A(n639), .Y(n1310) );
  AOI22X1 U1187 ( .A0(dR_reg[1]), .A1(n1352), .B0(deg_Ri[1]), .B1(n1316), .Y(
        n639) );
  INVX1 U1188 ( .A(n640), .Y(n1311) );
  AOI22X1 U1189 ( .A0(dR_reg[2]), .A1(n1357), .B0(deg_Ri[2]), .B1(n1315), .Y(
        n640) );
  INVX1 U1190 ( .A(n641), .Y(n1312) );
  AOI22X1 U1191 ( .A0(dR_reg[3]), .A1(n1360), .B0(deg_Ri[3]), .B1(n1316), .Y(
        n641) );
  INVX1 U1192 ( .A(n642), .Y(n1313) );
  AOI22X1 U1193 ( .A0(dR_reg[4]), .A1(n1362), .B0(deg_Ri[4]), .B1(n1046), .Y(
        n642) );
  INVX1 U1194 ( .A(n395), .Y(n1063) );
  AOI22X1 U1195 ( .A0(n1375), .A1(LLL2[4]), .B0(n1325), .B1(LLL1[4]), .Y(n395)
         );
  INVX1 U1196 ( .A(n405), .Y(n1073) );
  AOI22X1 U1197 ( .A0(n1378), .A1(LLL2[3]), .B0(n1325), .B1(LLL1[3]), .Y(n405)
         );
  INVX1 U1198 ( .A(n15), .Y(n682) );
  AOI22X1 U1199 ( .A0(n806), .A1(DR7[3]), .B0(DR8[3]), .B1(n1348), .Y(n15) );
  INVX1 U1200 ( .A(n23), .Y(n690) );
  AOI22X1 U1201 ( .A0(n806), .A1(DR7[2]), .B0(DR8[2]), .B1(n1342), .Y(n23) );
  INVX1 U1202 ( .A(n31), .Y(n698) );
  AOI22X1 U1203 ( .A0(n806), .A1(DR7[1]), .B0(DR8[1]), .B1(n1348), .Y(n31) );
  INVX1 U1204 ( .A(n39), .Y(n706) );
  AOI22X1 U1205 ( .A0(n806), .A1(DR7[0]), .B0(DR8[0]), .B1(n1344), .Y(n39) );
  INVX1 U1206 ( .A(n47), .Y(n714) );
  AOI22X1 U1207 ( .A0(n806), .A1(DQ7[4]), .B0(DQ8[4]), .B1(n1346), .Y(n47) );
  INVX1 U1208 ( .A(n55), .Y(n722) );
  AOI22X1 U1209 ( .A0(n814), .A1(DQ7[3]), .B0(DQ8[3]), .B1(n1352), .Y(n55) );
  INVX1 U1210 ( .A(n63), .Y(n730) );
  AOI22X1 U1211 ( .A0(n814), .A1(DQ7[2]), .B0(DQ8[2]), .B1(n1358), .Y(n63) );
  INVX1 U1212 ( .A(n71), .Y(n738) );
  AOI22X1 U1213 ( .A0(n814), .A1(DQ7[1]), .B0(DQ8[1]), .B1(n1366), .Y(n71) );
  INVX1 U1214 ( .A(n79), .Y(n746) );
  AOI22X1 U1215 ( .A0(n814), .A1(DQ7[0]), .B0(DQ8[0]), .B1(n1388), .Y(n79) );
  INVX1 U1216 ( .A(n87), .Y(n754) );
  AOI22X1 U1217 ( .A0(n814), .A1(ST1), .B0(ST2), .B1(n1369), .Y(n87) );
  INVX1 U1218 ( .A(n99), .Y(n767) );
  AOI22X1 U1219 ( .A0(n830), .A1(R7[12]), .B0(R8[12]), .B1(n1401), .Y(n99) );
  INVX1 U1220 ( .A(n107), .Y(n775) );
  AOI22X1 U1221 ( .A0(n838), .A1(R7[11]), .B0(R8[11]), .B1(n1377), .Y(n107) );
  INVX1 U1222 ( .A(n115), .Y(n783) );
  AOI22X1 U1223 ( .A0(n846), .A1(R7[10]), .B0(R8[10]), .B1(n1388), .Y(n115) );
  INVX1 U1224 ( .A(n123), .Y(n791) );
  AOI22X1 U1225 ( .A0(n846), .A1(R7[9]), .B0(R8[9]), .B1(n1382), .Y(n123) );
  INVX1 U1226 ( .A(n131), .Y(n799) );
  AOI22X1 U1227 ( .A0(n986), .A1(R7[8]), .B0(R8[8]), .B1(n1389), .Y(n131) );
  INVX1 U1228 ( .A(n139), .Y(n807) );
  AOI22X1 U1229 ( .A0(n994), .A1(R7[7]), .B0(R8[7]), .B1(n1389), .Y(n139) );
  INVX1 U1230 ( .A(n147), .Y(n815) );
  AOI22X1 U1231 ( .A0(n994), .A1(R7[6]), .B0(R8[6]), .B1(n1353), .Y(n147) );
  INVX1 U1232 ( .A(n155), .Y(n823) );
  AOI22X1 U1233 ( .A0(n996), .A1(R7[5]), .B0(R8[5]), .B1(n1342), .Y(n155) );
  INVX1 U1234 ( .A(n163), .Y(n831) );
  AOI22X1 U1235 ( .A0(n1004), .A1(R7[4]), .B0(R8[4]), .B1(n1404), .Y(n163) );
  INVX1 U1236 ( .A(n171), .Y(n839) );
  AOI22X1 U1237 ( .A0(n1016), .A1(R7[3]), .B0(R8[3]), .B1(n1382), .Y(n171) );
  INVX1 U1238 ( .A(n179), .Y(n847) );
  AOI22X1 U1239 ( .A0(n1026), .A1(R7[2]), .B0(R8[2]), .B1(n1401), .Y(n179) );
  INVX1 U1240 ( .A(n187), .Y(n855) );
  AOI22X1 U1241 ( .A0(n1024), .A1(R7[1]), .B0(R8[1]), .B1(n1337), .Y(n187) );
  INVX1 U1242 ( .A(n195), .Y(n863) );
  AOI22X1 U1243 ( .A0(n1014), .A1(R7[0]), .B0(R8[0]), .B1(n1400), .Y(n195) );
  INVX1 U1244 ( .A(n203), .Y(n871) );
  AOI22X1 U1245 ( .A0(n1026), .A1(Q7[12]), .B0(Q8[12]), .B1(n1403), .Y(n203)
         );
  INVX1 U1246 ( .A(n211), .Y(n879) );
  AOI22X1 U1247 ( .A0(n1024), .A1(Q7[11]), .B0(Q8[11]), .B1(n1379), .Y(n211)
         );
  INVX1 U1248 ( .A(n219), .Y(n887) );
  AOI22X1 U1249 ( .A0(n1006), .A1(Q7[10]), .B0(Q8[10]), .B1(n1359), .Y(n219)
         );
  INVX1 U1250 ( .A(n227), .Y(n895) );
  AOI22X1 U1251 ( .A0(n1004), .A1(Q7[9]), .B0(Q8[9]), .B1(n1408), .Y(n227) );
  INVX1 U1252 ( .A(n235), .Y(n903) );
  AOI22X1 U1253 ( .A0(n662), .A1(Q7[8]), .B0(Q8[8]), .B1(n1342), .Y(n235) );
  INVX1 U1254 ( .A(n243), .Y(n911) );
  AOI22X1 U1255 ( .A0(n661), .A1(Q7[7]), .B0(Q8[7]), .B1(n1368), .Y(n243) );
  INVX1 U1256 ( .A(n251), .Y(n919) );
  AOI22X1 U1257 ( .A0(n660), .A1(Q7[6]), .B0(Q8[6]), .B1(n1366), .Y(n251) );
  INVX1 U1258 ( .A(n259), .Y(n927) );
  AOI22X1 U1259 ( .A0(n660), .A1(Q7[5]), .B0(Q8[5]), .B1(n1365), .Y(n259) );
  INVX1 U1260 ( .A(n267), .Y(n935) );
  AOI22X1 U1261 ( .A0(n659), .A1(Q7[4]), .B0(Q8[4]), .B1(n1362), .Y(n267) );
  INVX1 U1262 ( .A(n275), .Y(n943) );
  AOI22X1 U1263 ( .A0(n658), .A1(Q7[3]), .B0(Q8[3]), .B1(n1359), .Y(n275) );
  INVX1 U1264 ( .A(n283), .Y(n951) );
  AOI22X1 U1265 ( .A0(n658), .A1(Q7[2]), .B0(Q8[2]), .B1(n1354), .Y(n283) );
  INVX1 U1266 ( .A(n291), .Y(n959) );
  AOI22X1 U1267 ( .A0(n657), .A1(Q7[1]), .B0(Q8[1]), .B1(n1351), .Y(n291) );
  INVX1 U1268 ( .A(n299), .Y(n967) );
  AOI22X1 U1269 ( .A0(n656), .A1(Q7[0]), .B0(Q8[0]), .B1(n1353), .Y(n299) );
  INVX1 U1270 ( .A(n309), .Y(n977) );
  AOI22X1 U1271 ( .A0(n655), .A1(LLL7[12]), .B0(LLL8[12]), .B1(n1345), .Y(n309) );
  INVX1 U1272 ( .A(n317), .Y(n985) );
  AOI22X1 U1273 ( .A0(n655), .A1(L1[11]), .B0(L2[11]), .B1(n1343), .Y(n317) );
  INVX1 U1274 ( .A(n319), .Y(n987) );
  AOI22X1 U1275 ( .A0(n655), .A1(LLL7[11]), .B0(LLL8[11]), .B1(n1343), .Y(n319) );
  INVX1 U1276 ( .A(n327), .Y(n995) );
  AOI22X1 U1277 ( .A0(n655), .A1(L1[10]), .B0(L2[10]), .B1(n1347), .Y(n327) );
  INVX1 U1278 ( .A(n329), .Y(n997) );
  AOI22X1 U1279 ( .A0(n655), .A1(LLL7[10]), .B0(LLL8[10]), .B1(n1342), .Y(n329) );
  INVX1 U1280 ( .A(n337), .Y(n1005) );
  AOI22X1 U1281 ( .A0(n655), .A1(L1[9]), .B0(L2[9]), .B1(n1345), .Y(n337) );
  INVX1 U1282 ( .A(n339), .Y(n1007) );
  AOI22X1 U1283 ( .A0(n655), .A1(LLL7[9]), .B0(LLL8[9]), .B1(n1341), .Y(n339)
         );
  INVX1 U1284 ( .A(n347), .Y(n1015) );
  AOI22X1 U1285 ( .A0(n653), .A1(L1[8]), .B0(L2[8]), .B1(n1404), .Y(n347) );
  INVX1 U1286 ( .A(n349), .Y(n1017) );
  AOI22X1 U1287 ( .A0(n653), .A1(LLL7[8]), .B0(LLL8[8]), .B1(n1400), .Y(n349)
         );
  INVX1 U1288 ( .A(n357), .Y(n1025) );
  AOI22X1 U1289 ( .A0(n653), .A1(L1[7]), .B0(L2[7]), .B1(n1353), .Y(n357) );
  INVX1 U1290 ( .A(n359), .Y(n1027) );
  AOI22X1 U1291 ( .A0(n653), .A1(LLL7[7]), .B0(LLL8[7]), .B1(n1344), .Y(n359)
         );
  INVX1 U1292 ( .A(n367), .Y(n1035) );
  AOI22X1 U1293 ( .A0(n653), .A1(L1[6]), .B0(L2[6]), .B1(n1347), .Y(n367) );
  INVX1 U1294 ( .A(n369), .Y(n1037) );
  AOI22X1 U1295 ( .A0(n653), .A1(LLL7[6]), .B0(LLL8[6]), .B1(n1349), .Y(n369)
         );
  INVX1 U1296 ( .A(n377), .Y(n1045) );
  AOI22X1 U1297 ( .A0(n653), .A1(L1[5]), .B0(L2[5]), .B1(n1356), .Y(n377) );
  INVX1 U1298 ( .A(n379), .Y(n1047) );
  AOI22X1 U1299 ( .A0(n653), .A1(LLL7[5]), .B0(LLL8[5]), .B1(n1355), .Y(n379)
         );
  INVX1 U1300 ( .A(n387), .Y(n1055) );
  AOI22X1 U1301 ( .A0(n652), .A1(L1[4]), .B0(L2[4]), .B1(n1361), .Y(n387) );
  INVX1 U1302 ( .A(n389), .Y(n1057) );
  AOI22X1 U1303 ( .A0(n652), .A1(LLL7[4]), .B0(LLL8[4]), .B1(n1361), .Y(n389)
         );
  INVX1 U1304 ( .A(n399), .Y(n1067) );
  AOI22X1 U1305 ( .A0(n652), .A1(LLL7[3]), .B0(LLL8[3]), .B1(n1351), .Y(n399)
         );
  INVX1 U1306 ( .A(n407), .Y(n1075) );
  AOI22X1 U1307 ( .A0(n652), .A1(L1[2]), .B0(L2[2]), .B1(n1350), .Y(n407) );
  INVX1 U1308 ( .A(n409), .Y(n1077) );
  AOI22X1 U1309 ( .A0(n652), .A1(LLL7[2]), .B0(LLL8[2]), .B1(n1349), .Y(n409)
         );
  INVX1 U1310 ( .A(n417), .Y(n1085) );
  AOI22X1 U1311 ( .A0(n652), .A1(L1[1]), .B0(L2[1]), .B1(n1352), .Y(n417) );
  INVX1 U1312 ( .A(n419), .Y(n1087) );
  AOI22X1 U1313 ( .A0(n650), .A1(LLL7[1]), .B0(LLL8[1]), .B1(n1354), .Y(n419)
         );
  INVX1 U1314 ( .A(n427), .Y(n1095) );
  AOI22X1 U1315 ( .A0(n650), .A1(L1[0]), .B0(L2[0]), .B1(n1360), .Y(n427) );
  INVX1 U1316 ( .A(n429), .Y(n1097) );
  AOI22X1 U1317 ( .A0(n650), .A1(LLL7[0]), .B0(LLL8[0]), .B1(n1359), .Y(n429)
         );
  INVX1 U1318 ( .A(n437), .Y(n1105) );
  AOI22X1 U1319 ( .A0(n650), .A1(U7[12]), .B0(U8[12]), .B1(n1364), .Y(n437) );
  INVX1 U1320 ( .A(n445), .Y(n1113) );
  AOI22X1 U1321 ( .A0(n649), .A1(Uout[12]), .B0(Uout_temp[12]), .B1(n1367), 
        .Y(n445) );
  INVX1 U1322 ( .A(n446), .Y(n1114) );
  AOI22X1 U1323 ( .A0(n649), .A1(U7[11]), .B0(U8[11]), .B1(n1368), .Y(n446) );
  INVX1 U1324 ( .A(n454), .Y(n1122) );
  AOI22X1 U1325 ( .A0(n806), .A1(Uout[11]), .B0(Uout_temp[11]), .B1(n1402), 
        .Y(n454) );
  INVX1 U1326 ( .A(n455), .Y(n1123) );
  AOI22X1 U1327 ( .A0(n798), .A1(U7[10]), .B0(U8[10]), .B1(n1356), .Y(n455) );
  INVX1 U1328 ( .A(n463), .Y(n1131) );
  AOI22X1 U1329 ( .A0(n798), .A1(Uout[10]), .B0(Uout_temp[10]), .B1(n1378), 
        .Y(n463) );
  INVX1 U1330 ( .A(n464), .Y(n1132) );
  AOI22X1 U1331 ( .A0(n798), .A1(U7[9]), .B0(U8[9]), .B1(n1376), .Y(n464) );
  INVX1 U1332 ( .A(n472), .Y(n1140) );
  AOI22X1 U1333 ( .A0(n790), .A1(Uout[9]), .B0(Uout_temp[9]), .B1(n1404), .Y(
        n472) );
  INVX1 U1334 ( .A(n473), .Y(n1141) );
  AOI22X1 U1335 ( .A0(n790), .A1(U7[8]), .B0(U8[8]), .B1(n1404), .Y(n473) );
  INVX1 U1336 ( .A(n481), .Y(n1149) );
  AOI22X1 U1337 ( .A0(n782), .A1(Uout[8]), .B0(Uout_temp[8]), .B1(n1401), .Y(
        n481) );
  INVX1 U1338 ( .A(n482), .Y(n1150) );
  AOI22X1 U1339 ( .A0(n782), .A1(U7[7]), .B0(U8[7]), .B1(n1389), .Y(n482) );
  INVX1 U1340 ( .A(n490), .Y(n1158) );
  AOI22X1 U1341 ( .A0(n670), .A1(Uout[7]), .B0(Uout_temp[7]), .B1(n1358), .Y(
        n490) );
  INVX1 U1342 ( .A(n491), .Y(n1159) );
  AOI22X1 U1343 ( .A0(n670), .A1(U7[6]), .B0(U8[6]), .B1(n1352), .Y(n491) );
  INVX1 U1344 ( .A(n499), .Y(n1167) );
  AOI22X1 U1345 ( .A0(n669), .A1(Uout[6]), .B0(Uout_temp[6]), .B1(n1352), .Y(
        n499) );
  INVX1 U1346 ( .A(n500), .Y(n1168) );
  AOI22X1 U1347 ( .A0(n669), .A1(U7[5]), .B0(U8[5]), .B1(n1388), .Y(n500) );
  INVX1 U1348 ( .A(n508), .Y(n1176) );
  AOI22X1 U1349 ( .A0(n668), .A1(Uout[5]), .B0(Uout_temp[5]), .B1(n1403), .Y(
        n508) );
  INVX1 U1350 ( .A(n509), .Y(n1177) );
  AOI22X1 U1351 ( .A0(n668), .A1(U7[4]), .B0(U8[4]), .B1(n1401), .Y(n509) );
  INVX1 U1352 ( .A(n517), .Y(n1185) );
  AOI22X1 U1353 ( .A0(n667), .A1(Uout[4]), .B0(Uout_temp[4]), .B1(n1403), .Y(
        n517) );
  INVX1 U1354 ( .A(n518), .Y(n1186) );
  AOI22X1 U1355 ( .A0(n667), .A1(U7[3]), .B0(U8[3]), .B1(n1402), .Y(n518) );
  INVX1 U1356 ( .A(n527), .Y(n1195) );
  AOI22X1 U1357 ( .A0(n666), .A1(U7[2]), .B0(U8[2]), .B1(n1359), .Y(n527) );
  INVX1 U1358 ( .A(n536), .Y(n1204) );
  AOI22X1 U1359 ( .A0(n665), .A1(U7[1]), .B0(U8[1]), .B1(n1403), .Y(n536) );
  INVX1 U1360 ( .A(n544), .Y(n1212) );
  AOI22X1 U1361 ( .A0(n665), .A1(Uout[1]), .B0(Uout_temp[1]), .B1(n1388), .Y(
        n544) );
  INVX1 U1362 ( .A(n545), .Y(n1213) );
  AOI22X1 U1363 ( .A0(n664), .A1(U7[0]), .B0(U8[0]), .B1(n1402), .Y(n545) );
  INVX1 U1364 ( .A(n553), .Y(n1221) );
  AOI22X1 U1365 ( .A0(n664), .A1(Uout[0]), .B0(Uout_temp[0]), .B1(n1378), .Y(
        n553) );
  INVX1 U1366 ( .A(n594), .Y(n1263) );
  AOI22X1 U1367 ( .A0(Lin[0]), .A1(n647), .B0(Lin_reg[0]), .B1(n1401), .Y(n594) );
  INVX1 U1368 ( .A(n595), .Y(n1264) );
  AOI22X1 U1369 ( .A0(Lin[1]), .A1(n647), .B0(Lin_reg[1]), .B1(n1355), .Y(n595) );
  INVX1 U1370 ( .A(n596), .Y(n1265) );
  AOI22X1 U1371 ( .A0(Lin[2]), .A1(n647), .B0(Lin_reg[2]), .B1(n1357), .Y(n596) );
  INVX1 U1372 ( .A(n597), .Y(n1266) );
  AOI22X1 U1373 ( .A0(Lin[3]), .A1(n647), .B0(Lin_reg[3]), .B1(n1362), .Y(n597) );
  INVX1 U1374 ( .A(n598), .Y(n1267) );
  AOI22X1 U1375 ( .A0(Lin[4]), .A1(n647), .B0(Lin_reg[4]), .B1(n1358), .Y(n598) );
  INVX1 U1376 ( .A(n599), .Y(n1268) );
  AOI22X1 U1377 ( .A0(Lin[5]), .A1(n647), .B0(Lin_reg[5]), .B1(n1360), .Y(n599) );
  INVX1 U1378 ( .A(n600), .Y(n1269) );
  AOI22X1 U1379 ( .A0(Lin[6]), .A1(n647), .B0(Lin_reg[6]), .B1(n1364), .Y(n600) );
  INVX1 U1380 ( .A(n601), .Y(n1270) );
  AOI22X1 U1381 ( .A0(Lin[7]), .A1(n647), .B0(Lin_reg[7]), .B1(n1363), .Y(n601) );
  INVX1 U1382 ( .A(n602), .Y(n1271) );
  AOI22X1 U1383 ( .A0(Lin[8]), .A1(n647), .B0(Lin_reg[8]), .B1(n1363), .Y(n602) );
  INVX1 U1384 ( .A(n603), .Y(n1272) );
  AOI22X1 U1385 ( .A0(Lin[9]), .A1(n646), .B0(Lin_reg[9]), .B1(n1367), .Y(n603) );
  INVX1 U1386 ( .A(n604), .Y(n1273) );
  AOI22X1 U1387 ( .A0(Lin[10]), .A1(n646), .B0(Lin_reg[10]), .B1(n1365), .Y(
        n604) );
  INVX1 U1388 ( .A(n605), .Y(n1274) );
  AOI22X1 U1389 ( .A0(Lin[11]), .A1(n647), .B0(Lin_reg[11]), .B1(n1369), .Y(
        n605) );
  INVX1 U1390 ( .A(n606), .Y(n1275) );
  AOI22X1 U1391 ( .A0(Lin[12]), .A1(n646), .B0(Lin_reg[12]), .B1(n1400), .Y(
        n606) );
  INVX1 U1392 ( .A(n560), .Y(n1229) );
  AOI22X1 U1393 ( .A0(n1339), .A1(START1), .B0(st_out), .B1(n1056), .Y(n560)
         );
  INVX1 U1394 ( .A(n89), .Y(n757) );
  AOI22X1 U1395 ( .A0(n814), .A1(s_reg[0]), .B0(n1386), .B1(s_reg[1]), .Y(n89)
         );
  INVX1 U1396 ( .A(n554), .Y(n1223) );
  AOI22X1 U1397 ( .A0(n664), .A1(START6), .B0(n1406), .B1(START7), .Y(n554) );
  INVX1 U1398 ( .A(n561), .Y(n1231) );
  AOI22X1 U1399 ( .A0(n662), .A1(stop3[0]), .B0(n1376), .B1(stop3[1]), .Y(n561) );
  INVX1 U1400 ( .A(n563), .Y(n1234) );
  AOI22X1 U1401 ( .A0(n668), .A1(stop2[0]), .B0(n1336), .B1(stop2[1]), .Y(n563) );
  INVX1 U1402 ( .A(n565), .Y(n1237) );
  AOI22X1 U1403 ( .A0(n650), .A1(stop1[0]), .B0(n1406), .B1(stop1[1]), .Y(n565) );
  INVX1 U1404 ( .A(N99), .Y(n1408) );
endmodule


module correct_module_4cells_p16 ( rstn, clk, start, gsynd, aadd1, aadd2, 
        aadd3, aadd4, aadd5, aadd6, aadd7, aadd8, sigma1, sigma2, sigma3, 
        sigma4, sigma5, sigma6, sigma7, sigma8, sigma9, sigma10, sigma11, 
        sigma12, sigma13, sigma14, sigma15, sigma16, err_count, pre_err, 
        error_occur, start_aadd, error_finish, error_number, e8, e_sum_r, 
        err_index, count, sig_all_zero, serr, Lout, enable_cs );
  input [12:0] gsynd;
  output [12:0] aadd1;
  output [12:0] aadd2;
  output [12:0] aadd3;
  output [12:0] aadd4;
  output [12:0] aadd5;
  output [12:0] aadd6;
  output [12:0] aadd7;
  output [12:0] aadd8;
  output [12:0] sigma1;
  output [12:0] sigma2;
  output [12:0] sigma3;
  output [12:0] sigma4;
  output [12:0] sigma5;
  output [12:0] sigma6;
  output [12:0] sigma7;
  output [12:0] sigma8;
  output [12:0] sigma9;
  output [12:0] sigma10;
  output [12:0] sigma11;
  output [12:0] sigma12;
  output [12:0] sigma13;
  output [12:0] sigma14;
  output [12:0] sigma15;
  output [12:0] sigma16;
  output [12:0] err_count;
  output [3:0] error_number;
  output [3:0] e_sum_r;
  output [15:0] err_index;
  output [9:0] count;
  output [3:0] serr;
  output [12:0] Lout;
  input rstn, clk, start;
  output pre_err, error_occur, start_aadd, error_finish, e8, sig_all_zero,
         enable_cs;
  wire   N256, N257, N258, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1675, n1676,
         stop_i, start_eu, sel_ch, N263, N264, N266, N270, N271, N272, N273,
         N274, N275, N276, N277, N278, N279, N327, N449, N661, N662, N663,
         N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N810,
         N811, N812, N813, N814, N815, N816, N817, N1141, N1190, n72, n77, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n96, n97, n98, n99, n100, n101, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n121, n122, n123,
         n124, n125, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n152, n153, n154, n155, n156, n157, n160, n165, n172,
         n175, n181, n182, n183, n184, n185, n186, n192, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n204, n206, n208, n210, n211,
         n212, n214, n225, n235, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n286, n287, n288, n289, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n515, n516, n517, n518, n519, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n736,
         n737, n738, n739, n740, n741, n742, n743, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, \add_587/carry[5] , \add_587/carry[6] ,
         \add_587/carry[7] , \add_587/carry[8] , \add_587/carry[9] ,
         \add_587/carry[10] , \add_587/carry[11] , \add_587/carry[12] , n807,
         n808, n809, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n825, n827, n828, n829, n830, n834, n837,
         n838, n839, n841, n842, n843, n845, n848, n850, n852, n854, n856,
         n857, n858, n859, n860, n861, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n934, n935, n936, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643;
  wire   [12:0] Rin;
  wire   [12:0] Uin;
  wire   [12:0] err_loc0;
  wire   [12:0] err_loc1;
  wire   [12:0] err_loc2;
  wire   [12:0] err_loc3;
  wire   [12:0] err_loc4;
  wire   [12:0] err_loc5;
  wire   [12:0] err_loc6;
  wire   [12:0] err_loc7;
  wire   [12:0] err_loc8;
  assign serr[0] = N256;
  assign serr[1] = N257;
  assign serr[2] = N258;
  assign N1190 = start;
  assign err_count[4] = \add_587/carry[5] ;

  euclidean_4cells euclidean ( .deg_Ri({1'b1, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .deg_Qi({1'b0, 1'b1, 1'b1, 1'b1, 1'b1}), .stop_i(stop_i), .Rin({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        Rin[0]}), .Qin(gsynd), .Lin({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Uin({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, Uin[0]}), .start(
        start_eu), .start_cnt(n972), .Lout(Lout), .clk(clk), .reset(rstn) );
  chien_search_p16_t8 chien ( .lambda0(err_loc0), .lambda1(err_loc1), 
        .lambda2(err_loc2), .lambda3(err_loc3), .lambda4(err_loc4), .lambda5(
        err_loc5), .lambda6(err_loc6), .lambda7(err_loc7), .lambda8(err_loc8), 
        .enable(enable_cs), .sigma1({sigma1[12:9], n1644, sigma1[7:6], n1645, 
        sigma1[4:0]}), .sigma2({sigma2[12:7], n1646, sigma2[5:0]}), .sigma3(
        sigma3), .sigma4(sigma4), .sigma5(sigma5), .sigma6(sigma6), .sigma7(
        sigma7), .sigma8(sigma8), .sigma9({sigma9[12:6], n1647, sigma9[4], 
        n1648, sigma9[2:0]}), .sigma10(sigma10), .sigma11({sigma11[12:7], 
        n1649, sigma11[5], n1650, n1651, n1652, n1653, sigma11[0]}), .sigma12(
        {sigma12[12:5], n1654, sigma12[3:0]}), .sigma13(sigma13), .sigma14({
        sigma14[12], n1655, sigma14[10:2], n1656, n1657}), .sigma15({
        sigma15[12:6], n1658, sigma15[4:0]}), .sigma16(sigma16), .sel(sel_ch), 
        .clk(clk), .reset(rstn) );
  correct_module_4cells_p16_DW01_inc_0 add_266 ( .A({count[9:6], n1675, n952, 
        count[3:0]}), .SUM({N279, N278, N277, N276, N275, N274, N273, N272, 
        N271, N270}) );
  DFFRHQX1 start_eu_reg ( .D(n751), .CK(clk), .RN(rstn), .Q(start_eu) );
  DFFRHQX1 \Uin_reg[0]  ( .D(n752), .CK(clk), .RN(rstn), .Q(Uin[0]) );
  DFFSX1 \aadd_reg[5][9]  ( .D(n694), .CK(clk), .SN(rstn), .Q(aadd6[9]), .QN(
        n570) );
  DFFSX1 \aadd_reg[5][8]  ( .D(n692), .CK(clk), .SN(rstn), .Q(aadd6[8]), .QN(
        n568) );
  DFFSX1 \aadd_reg[5][10]  ( .D(n691), .CK(clk), .SN(rstn), .Q(aadd6[10]), 
        .QN(n567) );
  DFFSX1 \aadd_reg[1][10]  ( .D(n655), .CK(clk), .SN(rstn), .Q(aadd2[10]), 
        .QN(n531) );
  DFFSX1 \aadd_reg[1][8]  ( .D(n654), .CK(clk), .SN(rstn), .Q(aadd2[8]), .QN(
        n530) );
  DFFSX1 \aadd_reg[1][9]  ( .D(n653), .CK(clk), .SN(rstn), .Q(aadd2[9]), .QN(
        n529) );
  DFFSX1 \aadd_reg[7][9]  ( .D(n629), .CK(clk), .SN(rstn), .Q(aadd8[9]), .QN(
        n505) );
  DFFSX1 \aadd_reg[7][8]  ( .D(n627), .CK(clk), .SN(rstn), .Q(aadd8[8]), .QN(
        n503) );
  DFFSX1 \aadd_reg[7][10]  ( .D(n626), .CK(clk), .SN(rstn), .Q(aadd8[10]), 
        .QN(n502) );
  DFFSX1 \aadd_reg[3][9]  ( .D(n616), .CK(clk), .SN(rstn), .Q(aadd4[9]), .QN(
        n492) );
  DFFSX1 \aadd_reg[3][8]  ( .D(n614), .CK(clk), .SN(rstn), .Q(aadd4[8]), .QN(
        n490) );
  DFFSX1 \aadd_reg[3][10]  ( .D(n613), .CK(clk), .SN(rstn), .Q(aadd4[10]), 
        .QN(n489) );
  DFFSX1 \aadd_reg[4][9]  ( .D(n681), .CK(clk), .SN(rstn), .Q(aadd5[9]), .QN(
        n557) );
  DFFSX1 \aadd_reg[4][8]  ( .D(n679), .CK(clk), .SN(rstn), .Q(aadd5[8]), .QN(
        n555) );
  DFFSX1 \aadd_reg[4][10]  ( .D(n678), .CK(clk), .SN(rstn), .Q(aadd5[10]), 
        .QN(n554) );
  DFFSX1 \aadd_reg[0][10]  ( .D(n642), .CK(clk), .SN(rstn), .Q(aadd1[10]), 
        .QN(n518) );
  DFFSX1 \aadd_reg[0][8]  ( .D(n641), .CK(clk), .SN(rstn), .Q(aadd1[8]), .QN(
        n517) );
  DFFSX1 \aadd_reg[0][9]  ( .D(n640), .CK(clk), .SN(rstn), .Q(aadd1[9]), .QN(
        n516) );
  DFFSX1 \aadd_reg[6][9]  ( .D(n707), .CK(clk), .SN(rstn), .Q(aadd7[9]), .QN(
        n583) );
  DFFSX1 \aadd_reg[6][8]  ( .D(n705), .CK(clk), .SN(rstn), .Q(aadd7[8]), .QN(
        n581) );
  DFFSX1 \aadd_reg[6][10]  ( .D(n704), .CK(clk), .SN(rstn), .Q(aadd7[10]), 
        .QN(n580) );
  DFFSX1 \aadd_reg[2][10]  ( .D(n668), .CK(clk), .SN(rstn), .Q(aadd3[10]), 
        .QN(n544) );
  DFFSX1 \aadd_reg[2][8]  ( .D(n667), .CK(clk), .SN(rstn), .Q(aadd3[8]), .QN(
        n543) );
  DFFSX1 \aadd_reg[2][9]  ( .D(n666), .CK(clk), .SN(rstn), .Q(aadd3[9]), .QN(
        n542) );
  DFFSX1 stop_i_reg ( .D(n750), .CK(clk), .SN(rstn), .Q(stop_i), .QN(n607) );
  DFFSX1 \Rin_reg[0]  ( .D(n749), .CK(clk), .SN(rstn), .Q(Rin[0]), .QN(n606)
         );
  DFFRHQX1 \err_loc0_reg[12]  ( .D(n1512), .CK(clk), .RN(rstn), .Q(
        err_loc0[12]) );
  DFFRHQX1 \err_loc0_reg[11]  ( .D(n1521), .CK(clk), .RN(rstn), .Q(
        err_loc0[11]) );
  DFFRHQX1 \err_loc0_reg[10]  ( .D(n1530), .CK(clk), .RN(rstn), .Q(
        err_loc0[10]) );
  DFFRHQX1 \err_loc0_reg[9]  ( .D(n1539), .CK(clk), .RN(rstn), .Q(err_loc0[9])
         );
  DFFRHQX1 \err_loc0_reg[8]  ( .D(n1548), .CK(clk), .RN(rstn), .Q(err_loc0[8])
         );
  DFFRHQX1 \err_loc0_reg[7]  ( .D(n1557), .CK(clk), .RN(rstn), .Q(err_loc0[7])
         );
  DFFRHQX1 \err_loc0_reg[6]  ( .D(n1566), .CK(clk), .RN(rstn), .Q(err_loc0[6])
         );
  DFFRHQX1 \err_loc0_reg[5]  ( .D(n1575), .CK(clk), .RN(rstn), .Q(err_loc0[5])
         );
  DFFRHQX1 \err_loc0_reg[4]  ( .D(n1584), .CK(clk), .RN(rstn), .Q(err_loc0[4])
         );
  DFFRHQX1 \err_loc0_reg[3]  ( .D(n1593), .CK(clk), .RN(rstn), .Q(err_loc0[3])
         );
  DFFRHQX1 \err_loc0_reg[2]  ( .D(n1602), .CK(clk), .RN(rstn), .Q(err_loc0[2])
         );
  DFFRHQX1 \err_loc0_reg[1]  ( .D(n1611), .CK(clk), .RN(rstn), .Q(err_loc0[1])
         );
  DFFRHQX1 \err_loc0_reg[0]  ( .D(n1620), .CK(clk), .RN(rstn), .Q(err_loc0[0])
         );
  DFFSX1 \aadd_reg[5][6]  ( .D(n699), .CK(clk), .SN(rstn), .Q(aadd6[6]), .QN(
        n575) );
  DFFSX1 \aadd_reg[5][4]  ( .D(n698), .CK(clk), .SN(rstn), .Q(aadd6[4]), .QN(
        n574) );
  DFFSX1 \aadd_reg[5][2]  ( .D(n697), .CK(clk), .SN(rstn), .Q(aadd6[2]), .QN(
        n573) );
  DFFSX1 \aadd_reg[5][0]  ( .D(n696), .CK(clk), .SN(rstn), .Q(aadd6[0]), .QN(
        n572) );
  DFFSX1 \aadd_reg[5][11]  ( .D(n695), .CK(clk), .SN(rstn), .Q(aadd6[11]), 
        .QN(n571) );
  DFFSX1 \aadd_reg[5][7]  ( .D(n693), .CK(clk), .SN(rstn), .Q(aadd6[7]), .QN(
        n569) );
  DFFSX1 \aadd_reg[5][12]  ( .D(n690), .CK(clk), .SN(rstn), .Q(aadd6[12]), 
        .QN(n566) );
  DFFSX1 \aadd_reg[5][1]  ( .D(n689), .CK(clk), .SN(rstn), .Q(aadd6[1]), .QN(
        n565) );
  DFFSX1 \aadd_reg[5][3]  ( .D(n688), .CK(clk), .SN(rstn), .Q(aadd6[3]), .QN(
        n564) );
  DFFSX1 \aadd_reg[5][5]  ( .D(n687), .CK(clk), .SN(rstn), .Q(aadd6[5]), .QN(
        n563) );
  DFFSX1 \aadd_reg[1][7]  ( .D(n660), .CK(clk), .SN(rstn), .Q(aadd2[7]), .QN(
        n536) );
  DFFSX1 \aadd_reg[1][5]  ( .D(n659), .CK(clk), .SN(rstn), .Q(aadd2[5]), .QN(
        n535) );
  DFFSX1 \aadd_reg[1][3]  ( .D(n658), .CK(clk), .SN(rstn), .Q(aadd2[3]), .QN(
        n534) );
  DFFSX1 \aadd_reg[1][1]  ( .D(n657), .CK(clk), .SN(rstn), .Q(aadd2[1]), .QN(
        n533) );
  DFFSX1 \aadd_reg[1][12]  ( .D(n656), .CK(clk), .SN(rstn), .Q(aadd2[12]), 
        .QN(n532) );
  DFFSX1 \aadd_reg[1][11]  ( .D(n652), .CK(clk), .SN(rstn), .Q(aadd2[11]), 
        .QN(n528) );
  DFFSX1 \aadd_reg[1][0]  ( .D(n651), .CK(clk), .SN(rstn), .Q(aadd2[0]), .QN(
        n527) );
  DFFSX1 \aadd_reg[1][2]  ( .D(n650), .CK(clk), .SN(rstn), .Q(aadd2[2]), .QN(
        n526) );
  DFFSX1 \aadd_reg[1][4]  ( .D(n649), .CK(clk), .SN(rstn), .Q(aadd2[4]), .QN(
        n525) );
  DFFSX1 \aadd_reg[1][6]  ( .D(n648), .CK(clk), .SN(rstn), .Q(aadd2[6]), .QN(
        n524) );
  DFFSX1 \aadd_reg[7][6]  ( .D(n634), .CK(clk), .SN(rstn), .Q(aadd8[6]), .QN(
        n510) );
  DFFSX1 \aadd_reg[7][4]  ( .D(n633), .CK(clk), .SN(rstn), .Q(aadd8[4]), .QN(
        n509) );
  DFFSX1 \aadd_reg[7][2]  ( .D(n632), .CK(clk), .SN(rstn), .Q(aadd8[2]), .QN(
        n508) );
  DFFSX1 \aadd_reg[7][0]  ( .D(n631), .CK(clk), .SN(rstn), .Q(aadd8[0]), .QN(
        n507) );
  DFFSX1 \aadd_reg[7][11]  ( .D(n630), .CK(clk), .SN(rstn), .Q(aadd8[11]), 
        .QN(n506) );
  DFFSX1 \aadd_reg[7][7]  ( .D(n628), .CK(clk), .SN(rstn), .Q(aadd8[7]), .QN(
        n504) );
  DFFSX1 \aadd_reg[7][12]  ( .D(n625), .CK(clk), .SN(rstn), .Q(aadd8[12]), 
        .QN(n501) );
  DFFSX1 \aadd_reg[7][1]  ( .D(n624), .CK(clk), .SN(rstn), .Q(aadd8[1]), .QN(
        n500) );
  DFFSX1 \aadd_reg[7][3]  ( .D(n623), .CK(clk), .SN(rstn), .Q(aadd8[3]), .QN(
        n499) );
  DFFSX1 \aadd_reg[7][5]  ( .D(n622), .CK(clk), .SN(rstn), .Q(aadd8[5]), .QN(
        n498) );
  DFFSX1 \aadd_reg[3][6]  ( .D(n621), .CK(clk), .SN(rstn), .Q(aadd4[6]), .QN(
        n497) );
  DFFSX1 \aadd_reg[3][4]  ( .D(n620), .CK(clk), .SN(rstn), .Q(aadd4[4]), .QN(
        n496) );
  DFFSX1 \aadd_reg[3][2]  ( .D(n619), .CK(clk), .SN(rstn), .Q(aadd4[2]), .QN(
        n495) );
  DFFSX1 \aadd_reg[3][0]  ( .D(n618), .CK(clk), .SN(rstn), .Q(aadd4[0]), .QN(
        n494) );
  DFFSX1 \aadd_reg[3][11]  ( .D(n617), .CK(clk), .SN(rstn), .Q(aadd4[11]), 
        .QN(n493) );
  DFFSX1 \aadd_reg[3][7]  ( .D(n615), .CK(clk), .SN(rstn), .Q(aadd4[7]), .QN(
        n491) );
  DFFSX1 \aadd_reg[3][12]  ( .D(n612), .CK(clk), .SN(rstn), .Q(aadd4[12]), 
        .QN(n488) );
  DFFSX1 \aadd_reg[3][1]  ( .D(n611), .CK(clk), .SN(rstn), .Q(aadd4[1]), .QN(
        n487) );
  DFFSX1 \aadd_reg[3][3]  ( .D(n610), .CK(clk), .SN(rstn), .Q(aadd4[3]), .QN(
        n486) );
  DFFSX1 \aadd_reg[3][5]  ( .D(n609), .CK(clk), .SN(rstn), .Q(aadd4[5]), .QN(
        n485) );
  DFFSX1 \aadd_reg[4][6]  ( .D(n686), .CK(clk), .SN(rstn), .Q(aadd5[6]), .QN(
        n562) );
  DFFSX1 \aadd_reg[4][4]  ( .D(n685), .CK(clk), .SN(rstn), .Q(aadd5[4]), .QN(
        n561) );
  DFFSX1 \aadd_reg[4][2]  ( .D(n684), .CK(clk), .SN(rstn), .Q(aadd5[2]), .QN(
        n560) );
  DFFSX1 \aadd_reg[4][0]  ( .D(n683), .CK(clk), .SN(rstn), .Q(aadd5[0]), .QN(
        n559) );
  DFFSX1 \aadd_reg[4][11]  ( .D(n682), .CK(clk), .SN(rstn), .Q(aadd5[11]), 
        .QN(n558) );
  DFFSX1 \aadd_reg[4][7]  ( .D(n680), .CK(clk), .SN(rstn), .Q(aadd5[7]), .QN(
        n556) );
  DFFSX1 \aadd_reg[4][12]  ( .D(n677), .CK(clk), .SN(rstn), .Q(aadd5[12]), 
        .QN(n553) );
  DFFSX1 \aadd_reg[4][1]  ( .D(n676), .CK(clk), .SN(rstn), .Q(aadd5[1]), .QN(
        n552) );
  DFFSX1 \aadd_reg[4][3]  ( .D(n675), .CK(clk), .SN(rstn), .Q(aadd5[3]), .QN(
        n551) );
  DFFSX1 \aadd_reg[4][5]  ( .D(n674), .CK(clk), .SN(rstn), .Q(aadd5[5]), .QN(
        n550) );
  DFFSX1 \aadd_reg[0][7]  ( .D(n647), .CK(clk), .SN(rstn), .Q(aadd1[7]), .QN(
        n523) );
  DFFSX1 \aadd_reg[0][5]  ( .D(n646), .CK(clk), .SN(rstn), .Q(aadd1[5]), .QN(
        n522) );
  DFFSX1 \aadd_reg[0][3]  ( .D(n645), .CK(clk), .SN(rstn), .Q(aadd1[3]) );
  DFFSX1 \aadd_reg[0][1]  ( .D(n644), .CK(clk), .SN(rstn), .Q(aadd1[1]) );
  DFFSX1 \aadd_reg[0][12]  ( .D(n643), .CK(clk), .SN(rstn), .Q(aadd1[12]), 
        .QN(n519) );
  DFFSX1 \aadd_reg[0][11]  ( .D(n639), .CK(clk), .SN(rstn), .Q(aadd1[11]), 
        .QN(n515) );
  DFFSX1 \aadd_reg[0][0]  ( .D(n638), .CK(clk), .SN(rstn), .Q(aadd1[0]) );
  DFFSX1 \aadd_reg[0][2]  ( .D(n637), .CK(clk), .SN(rstn), .Q(aadd1[2]) );
  DFFSX1 \aadd_reg[0][4]  ( .D(n636), .CK(clk), .SN(rstn), .Q(aadd1[4]), .QN(
        n512) );
  DFFSX1 \aadd_reg[0][6]  ( .D(n635), .CK(clk), .SN(rstn), .Q(aadd1[6]), .QN(
        n511) );
  DFFSX1 \aadd_reg[6][6]  ( .D(n712), .CK(clk), .SN(rstn), .Q(aadd7[6]), .QN(
        n588) );
  DFFSX1 \aadd_reg[6][4]  ( .D(n711), .CK(clk), .SN(rstn), .Q(aadd7[4]), .QN(
        n587) );
  DFFSX1 \aadd_reg[6][2]  ( .D(n710), .CK(clk), .SN(rstn), .Q(aadd7[2]), .QN(
        n586) );
  DFFSX1 \aadd_reg[6][0]  ( .D(n709), .CK(clk), .SN(rstn), .Q(aadd7[0]), .QN(
        n585) );
  DFFSX1 \aadd_reg[6][11]  ( .D(n708), .CK(clk), .SN(rstn), .Q(aadd7[11]), 
        .QN(n584) );
  DFFSX1 \aadd_reg[6][7]  ( .D(n706), .CK(clk), .SN(rstn), .Q(aadd7[7]), .QN(
        n582) );
  DFFSX1 \aadd_reg[6][12]  ( .D(n703), .CK(clk), .SN(rstn), .Q(aadd7[12]), 
        .QN(n579) );
  DFFSX1 \aadd_reg[6][1]  ( .D(n702), .CK(clk), .SN(rstn), .Q(aadd7[1]), .QN(
        n578) );
  DFFSX1 \aadd_reg[6][3]  ( .D(n701), .CK(clk), .SN(rstn), .Q(aadd7[3]), .QN(
        n577) );
  DFFSX1 \aadd_reg[6][5]  ( .D(n700), .CK(clk), .SN(rstn), .Q(aadd7[5]), .QN(
        n576) );
  DFFSX1 \aadd_reg[2][7]  ( .D(n673), .CK(clk), .SN(rstn), .Q(aadd3[7]), .QN(
        n549) );
  DFFSX1 \aadd_reg[2][5]  ( .D(n672), .CK(clk), .SN(rstn), .Q(aadd3[5]), .QN(
        n548) );
  DFFSX1 \aadd_reg[2][3]  ( .D(n671), .CK(clk), .SN(rstn), .Q(aadd3[3]), .QN(
        n547) );
  DFFSX1 \aadd_reg[2][1]  ( .D(n670), .CK(clk), .SN(rstn), .Q(aadd3[1]), .QN(
        n546) );
  DFFSX1 \aadd_reg[2][12]  ( .D(n669), .CK(clk), .SN(rstn), .Q(aadd3[12]), 
        .QN(n545) );
  DFFSX1 \aadd_reg[2][11]  ( .D(n665), .CK(clk), .SN(rstn), .Q(aadd3[11]), 
        .QN(n541) );
  DFFSX1 \aadd_reg[2][0]  ( .D(n664), .CK(clk), .SN(rstn), .Q(aadd3[0]), .QN(
        n540) );
  DFFSX1 \aadd_reg[2][2]  ( .D(n663), .CK(clk), .SN(rstn), .Q(aadd3[2]), .QN(
        n539) );
  DFFSX1 \aadd_reg[2][4]  ( .D(n662), .CK(clk), .SN(rstn), .Q(aadd3[4]), .QN(
        n538) );
  DFFSX1 \aadd_reg[2][6]  ( .D(n661), .CK(clk), .SN(rstn), .Q(aadd3[6]), .QN(
        n537) );
  DFFSX1 e13_reg ( .D(n740), .CK(clk), .SN(rstn), .Q(n814), .QN(n596) );
  DFFRHQX1 \count_reg[1]  ( .D(n761), .CK(clk), .RN(rstn), .Q(count[1]) );
  DFFRHQX1 \count_reg[2]  ( .D(n760), .CK(clk), .RN(rstn), .Q(count[2]) );
  DFFRHQX1 \count_reg[3]  ( .D(n759), .CK(clk), .RN(rstn), .Q(count[3]) );
  DFFRHQX1 \count_reg[4]  ( .D(n758), .CK(clk), .RN(rstn), .Q(count[4]) );
  DFFRHQX1 \count_reg[5]  ( .D(n757), .CK(clk), .RN(rstn), .Q(n1675) );
  DFFRHQX1 \count_reg[6]  ( .D(n756), .CK(clk), .RN(rstn), .Q(count[6]) );
  DFFRHQX1 \count_reg[7]  ( .D(n755), .CK(clk), .RN(rstn), .Q(count[7]) );
  DFFRHQX1 \count_reg[8]  ( .D(n754), .CK(clk), .RN(rstn), .Q(count[8]) );
  DFFRHQX1 start_aadd_reg ( .D(n748), .CK(clk), .RN(rstn), .Q(start_aadd) );
  DFFRHQX1 \err_loc3_reg[9]  ( .D(n1542), .CK(clk), .RN(rstn), .Q(err_loc3[9])
         );
  DFFRHQX1 \err_loc8_reg[7]  ( .D(n1565), .CK(clk), .RN(rstn), .Q(err_loc8[7])
         );
  DFFRHQX1 sel_ch_reg ( .D(N449), .CK(clk), .RN(rstn), .Q(sel_ch) );
  DFFRHQX1 \err_loc5_reg[12]  ( .D(n1517), .CK(clk), .RN(rstn), .Q(
        err_loc5[12]) );
  DFFRHQX1 \err_loc7_reg[11]  ( .D(n1528), .CK(clk), .RN(rstn), .Q(
        err_loc7[11]) );
  DFFRHQX1 \err_loc6_reg[10]  ( .D(n1536), .CK(clk), .RN(rstn), .Q(
        err_loc6[10]) );
  DFFRHQX1 \err_loc7_reg[10]  ( .D(n1537), .CK(clk), .RN(rstn), .Q(
        err_loc7[10]) );
  DFFRHQX1 \err_loc6_reg[5]  ( .D(n1581), .CK(clk), .RN(rstn), .Q(err_loc6[5])
         );
  DFFRHQX1 \err_loc3_reg[2]  ( .D(n1605), .CK(clk), .RN(rstn), .Q(err_loc3[2])
         );
  DFFRHQX1 \err_loc1_reg[12]  ( .D(n1513), .CK(clk), .RN(rstn), .Q(
        err_loc1[12]) );
  DFFRHQX1 \err_loc2_reg[12]  ( .D(n1514), .CK(clk), .RN(rstn), .Q(
        err_loc2[12]) );
  DFFRHQX1 \err_loc8_reg[11]  ( .D(n1529), .CK(clk), .RN(rstn), .Q(
        err_loc8[11]) );
  DFFRHQX1 \err_loc3_reg[10]  ( .D(n1533), .CK(clk), .RN(rstn), .Q(
        err_loc3[10]) );
  DFFRHQX1 \err_loc5_reg[10]  ( .D(n1535), .CK(clk), .RN(rstn), .Q(
        err_loc5[10]) );
  DFFRHQX1 \err_loc7_reg[6]  ( .D(n1573), .CK(clk), .RN(rstn), .Q(err_loc7[6])
         );
  DFFRHQX1 \err_loc1_reg[5]  ( .D(n1576), .CK(clk), .RN(rstn), .Q(err_loc1[5])
         );
  DFFRHQX1 \err_loc2_reg[4]  ( .D(n1586), .CK(clk), .RN(rstn), .Q(err_loc2[4])
         );
  DFFRHQX1 \err_loc2_reg[3]  ( .D(n1595), .CK(clk), .RN(rstn), .Q(err_loc2[3])
         );
  DFFRHQX1 \err_loc6_reg[2]  ( .D(n1608), .CK(clk), .RN(rstn), .Q(err_loc6[2])
         );
  DFFRHQX1 \err_loc1_reg[1]  ( .D(n1612), .CK(clk), .RN(rstn), .Q(err_loc1[1])
         );
  DFFRHQX1 \err_loc6_reg[0]  ( .D(n1626), .CK(clk), .RN(rstn), .Q(err_loc6[0])
         );
  DFFRHQX1 \err_loc6_reg[9]  ( .D(n1545), .CK(clk), .RN(rstn), .Q(err_loc6[9])
         );
  DFFRHQX1 \err_loc8_reg[10]  ( .D(n1538), .CK(clk), .RN(rstn), .Q(
        err_loc8[10]) );
  DFFRHQX1 \err_loc3_reg[7]  ( .D(n1560), .CK(clk), .RN(rstn), .Q(err_loc3[7])
         );
  DFFRHQX1 \err_loc3_reg[8]  ( .D(n1551), .CK(clk), .RN(rstn), .Q(err_loc3[8])
         );
  DFFRHQX1 \err_loc4_reg[7]  ( .D(n1561), .CK(clk), .RN(rstn), .Q(err_loc4[7])
         );
  DFFRHQX1 \err_loc3_reg[11]  ( .D(n1524), .CK(clk), .RN(rstn), .Q(
        err_loc3[11]) );
  DFFRHQX1 \err_loc8_reg[9]  ( .D(n1547), .CK(clk), .RN(rstn), .Q(err_loc8[9])
         );
  DFFRHQX1 \err_loc5_reg[8]  ( .D(n1553), .CK(clk), .RN(rstn), .Q(err_loc5[8])
         );
  DFFRHQX1 \err_loc8_reg[8]  ( .D(n1556), .CK(clk), .RN(rstn), .Q(err_loc8[8])
         );
  DFFRHQX1 \err_loc6_reg[7]  ( .D(n1563), .CK(clk), .RN(rstn), .Q(err_loc6[7])
         );
  DFFRHQX1 \err_loc3_reg[6]  ( .D(n1569), .CK(clk), .RN(rstn), .Q(err_loc3[6])
         );
  DFFRHQX1 \err_loc4_reg[6]  ( .D(n1570), .CK(clk), .RN(rstn), .Q(err_loc4[6])
         );
  DFFRHQX1 \err_loc3_reg[5]  ( .D(n1578), .CK(clk), .RN(rstn), .Q(err_loc3[5])
         );
  DFFRHQX1 \err_loc3_reg[4]  ( .D(n1587), .CK(clk), .RN(rstn), .Q(err_loc3[4])
         );
  DFFRHQX1 \err_loc1_reg[3]  ( .D(n1594), .CK(clk), .RN(rstn), .Q(err_loc1[3])
         );
  DFFRHQX1 \err_loc3_reg[1]  ( .D(n1614), .CK(clk), .RN(rstn), .Q(err_loc3[1])
         );
  DFFRHQX1 \err_loc6_reg[1]  ( .D(n1617), .CK(clk), .RN(rstn), .Q(err_loc6[1])
         );
  DFFRHQX1 \err_loc1_reg[0]  ( .D(n1621), .CK(clk), .RN(rstn), .Q(err_loc1[0])
         );
  DFFRHQX1 \err_loc3_reg[0]  ( .D(n1623), .CK(clk), .RN(rstn), .Q(err_loc3[0])
         );
  DFFRHQX1 \err_loc5_reg[11]  ( .D(n1526), .CK(clk), .RN(rstn), .Q(
        err_loc5[11]) );
  DFFRHQX1 \err_loc3_reg[3]  ( .D(n1596), .CK(clk), .RN(rstn), .Q(err_loc3[3])
         );
  DFFRHQX1 \err_loc5_reg[0]  ( .D(n1625), .CK(clk), .RN(rstn), .Q(err_loc5[0])
         );
  DFFRHQX1 \err_loc4_reg[11]  ( .D(n1525), .CK(clk), .RN(rstn), .Q(
        err_loc4[11]) );
  DFFRHQX1 \err_loc1_reg[10]  ( .D(n1531), .CK(clk), .RN(rstn), .Q(
        err_loc1[10]) );
  DFFRHQX1 \err_loc7_reg[8]  ( .D(n1555), .CK(clk), .RN(rstn), .Q(err_loc7[8])
         );
  DFFRHQX1 \err_loc1_reg[6]  ( .D(n1567), .CK(clk), .RN(rstn), .Q(err_loc1[6])
         );
  DFFRHQX1 \err_loc8_reg[2]  ( .D(n1610), .CK(clk), .RN(rstn), .Q(err_loc8[2])
         );
  DFFRHQX1 \err_loc8_reg[1]  ( .D(n1619), .CK(clk), .RN(rstn), .Q(err_loc8[1])
         );
  DFFRHQX1 \count_reg[9]  ( .D(n753), .CK(clk), .RN(rstn), .Q(count[9]) );
  DFFRHQX1 \count_reg[0]  ( .D(n762), .CK(clk), .RN(rstn), .Q(count[0]) );
  DFFRHQX1 \err_loc6_reg[6]  ( .D(n1572), .CK(clk), .RN(rstn), .Q(err_loc6[6])
         );
  DFFRHQX1 \err_loc8_reg[5]  ( .D(n1583), .CK(clk), .RN(rstn), .Q(err_loc8[5])
         );
  DFFRHQX1 \err_loc1_reg[9]  ( .D(n1540), .CK(clk), .RN(rstn), .Q(err_loc1[9])
         );
  DFFRHQX1 \err_loc7_reg[9]  ( .D(n1546), .CK(clk), .RN(rstn), .Q(err_loc7[9])
         );
  DFFRHQX1 \err_loc2_reg[5]  ( .D(n1577), .CK(clk), .RN(rstn), .Q(err_loc2[5])
         );
  DFFRHQX1 \err_loc2_reg[0]  ( .D(n1622), .CK(clk), .RN(rstn), .Q(err_loc2[0])
         );
  DFFRHQX1 \err_loc4_reg[12]  ( .D(n1516), .CK(clk), .RN(rstn), .Q(
        err_loc4[12]) );
  DFFRHQX1 \err_loc5_reg[9]  ( .D(n1544), .CK(clk), .RN(rstn), .Q(err_loc5[9])
         );
  DFFRHQX1 \err_loc5_reg[7]  ( .D(n1562), .CK(clk), .RN(rstn), .Q(err_loc5[7])
         );
  DFFRHQX1 \err_loc7_reg[3]  ( .D(n1600), .CK(clk), .RN(rstn), .Q(err_loc7[3])
         );
  DFFRHQX1 \err_loc8_reg[3]  ( .D(n1601), .CK(clk), .RN(rstn), .Q(err_loc8[3])
         );
  DFFRHQX1 \err_loc2_reg[10]  ( .D(n1532), .CK(clk), .RN(rstn), .Q(
        err_loc2[10]) );
  DFFRHQX1 \err_loc4_reg[10]  ( .D(n1534), .CK(clk), .RN(rstn), .Q(
        err_loc4[10]) );
  DFFRHQX1 \err_loc6_reg[8]  ( .D(n1554), .CK(clk), .RN(rstn), .Q(err_loc6[8])
         );
  DFFRHQX1 \err_loc8_reg[4]  ( .D(n1592), .CK(clk), .RN(rstn), .Q(err_loc8[4])
         );
  DFFRHQX1 \err_loc4_reg[3]  ( .D(n1597), .CK(clk), .RN(rstn), .Q(err_loc4[3])
         );
  DFFRHQX1 \err_loc5_reg[3]  ( .D(n1598), .CK(clk), .RN(rstn), .Q(err_loc5[3])
         );
  DFFRHQX1 \err_loc8_reg[0]  ( .D(n1628), .CK(clk), .RN(rstn), .Q(err_loc8[0])
         );
  DFFRHQX1 \err_loc7_reg[2]  ( .D(n1609), .CK(clk), .RN(rstn), .Q(err_loc7[2])
         );
  DFFRHQX1 \err_loc8_reg[12]  ( .D(n1520), .CK(clk), .RN(rstn), .Q(
        err_loc8[12]) );
  DFFRHQX1 \err_loc6_reg[3]  ( .D(n1599), .CK(clk), .RN(rstn), .Q(err_loc6[3])
         );
  DFFRHQX1 \err_loc5_reg[1]  ( .D(n1616), .CK(clk), .RN(rstn), .Q(err_loc5[1])
         );
  DFFRHQX1 \err_loc2_reg[11]  ( .D(n1523), .CK(clk), .RN(rstn), .Q(
        err_loc2[11]) );
  DFFRHQX1 \err_loc6_reg[11]  ( .D(n1527), .CK(clk), .RN(rstn), .Q(
        err_loc6[11]) );
  DFFRHQX1 \err_loc1_reg[8]  ( .D(n1549), .CK(clk), .RN(rstn), .Q(err_loc1[8])
         );
  DFFRHQX1 \err_loc4_reg[8]  ( .D(n1552), .CK(clk), .RN(rstn), .Q(err_loc4[8])
         );
  DFFRHQX1 \err_loc1_reg[7]  ( .D(n1558), .CK(clk), .RN(rstn), .Q(err_loc1[7])
         );
  DFFRHQX1 \err_loc2_reg[7]  ( .D(n1559), .CK(clk), .RN(rstn), .Q(err_loc2[7])
         );
  DFFRHQX1 \err_loc7_reg[7]  ( .D(n1564), .CK(clk), .RN(rstn), .Q(err_loc7[7])
         );
  DFFRHQX1 \err_loc4_reg[5]  ( .D(n1579), .CK(clk), .RN(rstn), .Q(err_loc4[5])
         );
  DFFRHQX1 \err_loc1_reg[4]  ( .D(n1585), .CK(clk), .RN(rstn), .Q(err_loc1[4])
         );
  DFFRHQX1 \err_loc4_reg[4]  ( .D(n1588), .CK(clk), .RN(rstn), .Q(err_loc4[4])
         );
  DFFRHQX1 \err_loc1_reg[2]  ( .D(n1603), .CK(clk), .RN(rstn), .Q(err_loc1[2])
         );
  DFFRHQX1 \err_loc2_reg[2]  ( .D(n1604), .CK(clk), .RN(rstn), .Q(err_loc2[2])
         );
  DFFRHQX1 \err_loc5_reg[2]  ( .D(n1607), .CK(clk), .RN(rstn), .Q(err_loc5[2])
         );
  DFFRHQX1 \err_loc4_reg[1]  ( .D(n1615), .CK(clk), .RN(rstn), .Q(err_loc4[1])
         );
  DFFRHQX1 \err_loc4_reg[0]  ( .D(n1624), .CK(clk), .RN(rstn), .Q(err_loc4[0])
         );
  DFFRHQX1 \err_loc2_reg[9]  ( .D(n1541), .CK(clk), .RN(rstn), .Q(err_loc2[9])
         );
  DFFRHQX1 \err_loc4_reg[9]  ( .D(n1543), .CK(clk), .RN(rstn), .Q(err_loc4[9])
         );
  DFFRHQX1 \err_loc2_reg[6]  ( .D(n1568), .CK(clk), .RN(rstn), .Q(err_loc2[6])
         );
  DFFRHQX1 \err_loc5_reg[6]  ( .D(n1571), .CK(clk), .RN(rstn), .Q(err_loc5[6])
         );
  DFFRHQX1 \err_loc4_reg[2]  ( .D(n1606), .CK(clk), .RN(rstn), .Q(err_loc4[2])
         );
  DFFRHQX1 \err_loc5_reg[5]  ( .D(n1580), .CK(clk), .RN(rstn), .Q(err_loc5[5])
         );
  DFFRHQX1 \err_loc2_reg[8]  ( .D(n1550), .CK(clk), .RN(rstn), .Q(err_loc2[8])
         );
  DFFRHQX1 \err_loc1_reg[11]  ( .D(n1522), .CK(clk), .RN(rstn), .Q(
        err_loc1[11]) );
  DFFRHQX1 \err_loc7_reg[5]  ( .D(n1582), .CK(clk), .RN(rstn), .Q(err_loc7[5])
         );
  DFFRHQX1 \err_loc5_reg[4]  ( .D(n1589), .CK(clk), .RN(rstn), .Q(err_loc5[4])
         );
  DFFRHQX1 \err_loc2_reg[1]  ( .D(n1613), .CK(clk), .RN(rstn), .Q(err_loc2[1])
         );
  DFFRHQX1 \err_loc7_reg[1]  ( .D(n1618), .CK(clk), .RN(rstn), .Q(err_loc7[1])
         );
  DFFRHQX1 \err_loc7_reg[12]  ( .D(n1519), .CK(clk), .RN(rstn), .Q(
        err_loc7[12]) );
  DFFRHQX1 \err_loc8_reg[6]  ( .D(n1574), .CK(clk), .RN(rstn), .Q(err_loc8[6])
         );
  DFFRHQX1 \err_loc6_reg[4]  ( .D(n1590), .CK(clk), .RN(rstn), .Q(err_loc6[4])
         );
  DFFRHQX1 \err_loc7_reg[0]  ( .D(n1627), .CK(clk), .RN(rstn), .Q(err_loc7[0])
         );
  DFFRHQX1 \err_loc3_reg[12]  ( .D(n1515), .CK(clk), .RN(rstn), .Q(
        err_loc3[12]) );
  DFFSX1 \err_count_reg[5]  ( .D(n730), .CK(clk), .SN(rstn), .Q(err_count[5]), 
        .QN(n591) );
  DFFSX1 \err_count_reg[6]  ( .D(n729), .CK(clk), .SN(rstn), .Q(err_count[6]), 
        .QN(n590) );
  DFFSX1 \err_count_reg[4]  ( .D(n731), .CK(clk), .SN(rstn), .Q(
        \add_587/carry[5] ), .QN(n592) );
  DFFSX1 \err_count_reg[12]  ( .D(n723), .CK(clk), .SN(rstn), .Q(err_count[12]), .QN(n589) );
  DFFSX1 e9_reg ( .D(N1141), .CK(clk), .SN(rstn), .QN(n765) );
  DFFSX1 e14_reg ( .D(n739), .CK(clk), .SN(rstn), .Q(n822), .QN(n595) );
  DFFSX1 e6_reg ( .D(n717), .CK(clk), .SN(rstn), .Q(n815), .QN(n603) );
  DFFSX1 e10_reg ( .D(n743), .CK(clk), .SN(rstn), .Q(n900), .QN(n605) );
  DFFSX1 e7_reg ( .D(n716), .CK(clk), .SN(rstn), .Q(n899), .QN(n604) );
  DFFSX1 e8_reg ( .D(n715), .CK(clk), .SN(rstn), .Q(e8), .QN(n764) );
  DFFSX1 e16_reg ( .D(n608), .CK(clk), .SN(rstn), .QN(n593) );
  DFFRHQXL \e_sum_r_reg[2]  ( .D(n1509), .CK(clk), .RN(rstn), .Q(e_sum_r[2])
         );
  DFFSX1 e12_reg ( .D(n741), .CK(clk), .SN(rstn), .Q(n807), .QN(n597) );
  DFFRHQX1 \e_sum_r_reg[3]  ( .D(n1508), .CK(clk), .RN(rstn), .Q(e_sum_r[3])
         );
  DFFSX1 e15_reg ( .D(n738), .CK(clk), .SN(rstn), .Q(n821), .QN(n594) );
  DFFSX1 e11_reg ( .D(n742), .CK(clk), .SN(rstn), .Q(n820), .QN(n598) );
  DFFRHQX1 \e_sum_r_reg[1]  ( .D(n1510), .CK(clk), .RN(rstn), .Q(e_sum_r[1])
         );
  DFFRHQX1 \error_number_reg[3]  ( .D(n736), .CK(clk), .RN(rstn), .Q(
        error_number[3]) );
  DFFRHQX1 \err_loc7_reg[4]  ( .D(n1591), .CK(clk), .RN(rstn), .Q(err_loc7[4])
         );
  DFFRHQX1 \err_loc6_reg[12]  ( .D(n1518), .CK(clk), .RN(rstn), .Q(
        err_loc6[12]) );
  DFFSX1 e5_reg ( .D(n718), .CK(clk), .SN(rstn), .Q(n816), .QN(n599) );
  DFFRHQXL \e_sum_r_reg[0]  ( .D(n1511), .CK(clk), .RN(rstn), .Q(e_sum_r[0])
         );
  DFFRHQX2 \error_number_reg[2]  ( .D(n713), .CK(clk), .RN(rstn), .Q(N258) );
  DFFRHQX2 \err_count_reg[9]  ( .D(n726), .CK(clk), .RN(rstn), .Q(err_count[9]) );
  DFFRHQX2 \err_count_reg[11]  ( .D(n724), .CK(clk), .RN(rstn), .Q(
        err_count[11]) );
  DFFRHQX2 \err_count_reg[7]  ( .D(n728), .CK(clk), .RN(rstn), .Q(err_count[7]) );
  DFFRHQX2 \err_count_reg[10]  ( .D(n725), .CK(clk), .RN(rstn), .Q(
        err_count[10]) );
  DFFRHQX2 \err_count_reg[8]  ( .D(n727), .CK(clk), .RN(rstn), .Q(err_count[8]) );
  DFFRHQX1 \error_number_reg[1]  ( .D(n714), .CK(clk), .RN(rstn), .Q(N257) );
  DFFSX4 e3_reg ( .D(n720), .CK(clk), .SN(rstn), .Q(n809), .QN(n601) );
  DFFSX4 e1_reg ( .D(n722), .CK(clk), .SN(rstn), .Q(n813), .QN(n763) );
  DFFRHQX1 \error_number_reg[0]  ( .D(n737), .CK(clk), .RN(rstn), .Q(N256) );
  DFFSX1 e4_reg ( .D(n719), .CK(clk), .SN(rstn), .Q(n1506), .QN(n600) );
  DFFSX2 e2_reg ( .D(n721), .CK(clk), .SN(rstn), .Q(n823), .QN(n602) );
  INVX1 U763 ( .A(1'b0), .Y(err_index[0]) );
  INVX1 U765 ( .A(1'b0), .Y(err_index[1]) );
  INVX1 U767 ( .A(1'b0), .Y(err_index[2]) );
  INVX1 U769 ( .A(1'b0), .Y(err_index[3]) );
  INVX1 U771 ( .A(1'b0), .Y(err_index[4]) );
  INVX1 U773 ( .A(1'b0), .Y(err_index[5]) );
  INVX1 U775 ( .A(1'b0), .Y(err_index[6]) );
  INVX1 U777 ( .A(1'b0), .Y(err_index[7]) );
  INVX1 U779 ( .A(1'b0), .Y(err_index[8]) );
  INVX1 U781 ( .A(1'b0), .Y(err_index[9]) );
  INVX1 U783 ( .A(1'b0), .Y(err_index[10]) );
  INVX1 U785 ( .A(1'b0), .Y(err_index[11]) );
  INVX1 U787 ( .A(1'b0), .Y(err_index[12]) );
  INVX1 U789 ( .A(1'b0), .Y(err_index[13]) );
  INVX1 U791 ( .A(1'b0), .Y(err_index[14]) );
  INVX1 U793 ( .A(1'b0), .Y(err_index[15]) );
  INVX1 U795 ( .A(1'b1), .Y(err_count[0]) );
  INVX1 U797 ( .A(1'b1), .Y(err_count[1]) );
  INVX1 U799 ( .A(1'b1), .Y(err_count[2]) );
  INVX1 U801 ( .A(1'b1), .Y(err_count[3]) );
  NOR3XL U803 ( .A(n980), .B(n981), .C(1'b0), .Y(n979) );
  NAND2BXL U805 ( .AN(n1427), .B(n940), .Y(n1444) );
  INVX4 U806 ( .A(sig_all_zero), .Y(n1393) );
  AND4X4 U807 ( .A(n1121), .B(n883), .C(n1118), .D(n885), .Y(n850) );
  NOR4X1 U808 ( .A(sigma5[2]), .B(sigma5[3]), .C(sigma5[0]), .D(sigma5[1]), 
        .Y(n1080) );
  OAI2BB1X1 U809 ( .A0N(n1323), .A1N(n1320), .B0(n1316), .Y(n1378) );
  NAND2X2 U810 ( .A(n944), .B(n943), .Y(n1425) );
  INVX1 U811 ( .A(n1414), .Y(n1374) );
  INVX1 U812 ( .A(n1415), .Y(n1376) );
  NAND3X1 U813 ( .A(n1068), .B(n1067), .C(n1066), .Y(n1116) );
  NAND2X1 U814 ( .A(n1107), .B(n1106), .Y(n1392) );
  NOR3X1 U815 ( .A(sigma10[9]), .B(sigma10[7]), .C(sigma10[8]), .Y(n1001) );
  NOR3X1 U816 ( .A(sigma6[12]), .B(sigma6[10]), .C(sigma6[11]), .Y(n1069) );
  AND2X2 U817 ( .A(n1384), .B(n1394), .Y(n1347) );
  NAND2X1 U818 ( .A(n765), .B(n874), .Y(n1320) );
  OAI21X1 U819 ( .A0(n1412), .A1(n1411), .B0(n1413), .Y(n943) );
  NOR2X1 U820 ( .A(n971), .B(n1309), .Y(n856) );
  AND4X2 U821 ( .A(n199), .B(n820), .C(n807), .D(n142), .Y(n225) );
  INVX1 U822 ( .A(n204), .Y(n142) );
  OAI2BB1X2 U823 ( .A0N(n1390), .A1N(n1389), .B0(n1423), .Y(n1471) );
  OAI2BB1X1 U824 ( .A0N(n1356), .A1N(n1357), .B0(n1427), .Y(n1358) );
  NAND2X1 U825 ( .A(n1453), .B(n1471), .Y(n1454) );
  OR4X2 U826 ( .A(n1113), .B(n1280), .C(sigma15[11]), .D(sigma15[12]), .Y(
        n1114) );
  AOI21X1 U827 ( .A0(n808), .A1(n1633), .B0(n965), .Y(n902) );
  INVX1 U828 ( .A(count[9]), .Y(n808) );
  AOI2BB2X1 U829 ( .B0(n599), .B1(n1160), .A0N(n1327), .A1N(n857), .Y(n718) );
  NOR3X1 U830 ( .A(sigma11[11]), .B(n1301), .C(n1302), .Y(n817) );
  AND4X2 U831 ( .A(n987), .B(n986), .C(n989), .D(n988), .Y(n1121) );
  NAND3X1 U832 ( .A(e8), .B(n899), .C(n210), .Y(n204) );
  MX2X1 U833 ( .A(n901), .B(e_sum_r[1]), .S0(n971), .Y(n1510) );
  MX2X1 U834 ( .A(err_loc6[0]), .B(err_loc7[0]), .S0(n965), .Y(n1627) );
  NAND2BXL U835 ( .AN(n1130), .B(n1345), .Y(n1323) );
  XOR3X2 U836 ( .A(n1411), .B(n1414), .C(n1415), .Y(n1433) );
  NAND2XL U837 ( .A(n1340), .B(sig_all_zero), .Y(n875) );
  AOI2BB2X1 U838 ( .B0(n594), .B1(n1283), .A0N(n1282), .A1N(n1281), .Y(n738)
         );
  MX2X1 U839 ( .A(err_loc6[1]), .B(err_loc7[1]), .S0(n965), .Y(n1618) );
  NAND2BX1 U840 ( .AN(err_count[10]), .B(n978), .Y(n981) );
  AND2X2 U841 ( .A(n1387), .B(n1407), .Y(n1351) );
  NAND2X1 U842 ( .A(n1373), .B(n1372), .Y(n1379) );
  NAND2BX1 U843 ( .AN(n1369), .B(n1434), .Y(n1436) );
  NAND4X1 U844 ( .A(n809), .B(n813), .C(n600), .D(n823), .Y(n147) );
  NAND3X1 U845 ( .A(n974), .B(n1496), .C(n1497), .Y(n1487) );
  CLKINVX3 U846 ( .A(n1338), .Y(n1340) );
  OAI2BB1X1 U847 ( .A0N(n146), .A1N(n1309), .B0(n968), .Y(n1299) );
  MX2X1 U848 ( .A(err_loc7[0]), .B(err_loc8[0]), .S0(n965), .Y(n1628) );
  OAI2BB1X2 U849 ( .A0N(n599), .A1N(n1346), .B0(n1391), .Y(n1400) );
  OR4X2 U850 ( .A(n1140), .B(n1287), .C(n1655), .D(sigma14[12]), .Y(n1141) );
  NAND2XL U851 ( .A(n590), .B(n898), .Y(n984) );
  XOR2X1 U852 ( .A(n1457), .B(n1458), .Y(n1467) );
  NAND3XL U853 ( .A(n1480), .B(n1483), .C(n1445), .Y(n1446) );
  AOI2BB1X1 U854 ( .A0N(n266), .A1N(n267), .B0(n969), .Y(n950) );
  OAI2BB1X1 U855 ( .A0N(n77), .A1N(n875), .B0(n968), .Y(n1155) );
  MX2X1 U856 ( .A(err_loc1[0]), .B(err_loc2[0]), .S0(n965), .Y(n1622) );
  NAND2X1 U857 ( .A(n592), .B(n898), .Y(n982) );
  NAND4X1 U858 ( .A(n1057), .B(n1056), .C(n1055), .D(n1054), .Y(n818) );
  NAND2X1 U859 ( .A(n1387), .B(n1407), .Y(n889) );
  NAND2X1 U860 ( .A(n1377), .B(n1373), .Y(n1431) );
  AOI22XL U861 ( .A0(n127), .A1(err_count[9]), .B0(n128), .B1(N664), .Y(n89)
         );
  NOR3XL U862 ( .A(n206), .B(n593), .C(n594), .Y(n269) );
  NAND2BX1 U863 ( .AN(n1439), .B(n1442), .Y(n1450) );
  AOI2BB2X1 U864 ( .B0(n764), .B1(n1157), .A0N(n1312), .A1N(n857), .Y(n715) );
  MX2X1 U865 ( .A(err_loc7[1]), .B(err_loc8[1]), .S0(n965), .Y(n1619) );
  NAND4BXL U866 ( .AN(n1274), .B(n255), .C(n861), .D(n256), .Y(n1275) );
  OR2X2 U867 ( .A(n1117), .B(n1116), .Y(n819) );
  OAI2BB1X1 U868 ( .A0N(n599), .A1N(n1346), .B0(n1391), .Y(n812) );
  NAND2BX1 U869 ( .AN(n1380), .B(n1473), .Y(n945) );
  NAND2X1 U870 ( .A(n1033), .B(n1032), .Y(n1125) );
  NAND2X1 U871 ( .A(n591), .B(n592), .Y(\add_587/carry[6] ) );
  INVX1 U872 ( .A(n896), .Y(n128) );
  NAND3BXL U873 ( .AN(n1455), .B(n1440), .C(n1439), .Y(n1451) );
  AOI2BB1X1 U874 ( .A0N(n1284), .A1N(n822), .B0(n1290), .Y(n739) );
  MX2X1 U875 ( .A(err_loc0[0]), .B(err_loc1[0]), .S0(n965), .Y(n1621) );
  MX2X1 U876 ( .A(err_loc7[7]), .B(err_loc8[7]), .S0(n966), .Y(n1565) );
  CLKBUFXL U877 ( .A(n1658), .Y(sigma15[5]) );
  NOR2XL U878 ( .A(n1483), .B(n1482), .Y(n1484) );
  MXI2X1 U879 ( .A(n595), .B(n1142), .S0(n842), .Y(n1324) );
  INVX1 U880 ( .A(n1483), .Y(n811) );
  NAND3XL U881 ( .A(n1471), .B(n1470), .C(n1469), .Y(n1489) );
  OAI2BB1X2 U882 ( .A0N(n1479), .A1N(n1478), .B0(n1477), .Y(n1503) );
  NAND4X2 U883 ( .A(n1053), .B(n1052), .C(n1051), .D(n1050), .Y(n1058) );
  NAND2X1 U884 ( .A(n1318), .B(n1317), .Y(n1316) );
  CLKINVX3 U885 ( .A(n869), .Y(n870) );
  NAND2X1 U886 ( .A(n1315), .B(n1319), .Y(n1371) );
  OAI21X2 U887 ( .A0(n1326), .A1(n1325), .B0(n1324), .Y(n1373) );
  XOR3X2 U888 ( .A(n1410), .B(n828), .C(n827), .Y(n1412) );
  INVX1 U889 ( .A(n1409), .Y(n827) );
  NAND2X1 U890 ( .A(n1403), .B(n1404), .Y(n1410) );
  NAND2X1 U891 ( .A(sig_all_zero), .B(n1333), .Y(n1394) );
  CLKINVX3 U892 ( .A(n1411), .Y(n1402) );
  NAND2X2 U893 ( .A(n1425), .B(n1424), .Y(n1469) );
  INVXL U894 ( .A(n1366), .Y(n838) );
  OAI21XL U895 ( .A0(n1500), .A1(n1499), .B0(n1498), .Y(n1501) );
  NOR3X4 U896 ( .A(sigma9[10]), .B(sigma9[9]), .C(sigma9[12]), .Y(n869) );
  NAND4X2 U897 ( .A(n1003), .B(n1002), .C(n1001), .D(n1000), .Y(n1305) );
  NAND2X1 U898 ( .A(n1427), .B(n1426), .Y(n1491) );
  NOR3X1 U899 ( .A(n1049), .B(n1048), .C(n1047), .Y(n1102) );
  NOR2X2 U900 ( .A(n1105), .B(n1104), .Y(n1095) );
  NOR3X2 U901 ( .A(n1124), .B(n1133), .C(n1132), .Y(n1036) );
  INVX4 U902 ( .A(n874), .Y(n842) );
  NOR3X2 U903 ( .A(n602), .B(n601), .C(n763), .Y(n208) );
  NAND2BX2 U904 ( .AN(n1327), .B(n1345), .Y(n1391) );
  NAND2X1 U905 ( .A(n872), .B(n600), .Y(n1384) );
  NAND2XL U906 ( .A(n1676), .B(sig_all_zero), .Y(n872) );
  INVX1 U907 ( .A(n880), .Y(n881) );
  NAND4X1 U908 ( .A(n1013), .B(n1012), .C(n1011), .D(n1010), .Y(n1124) );
  NAND2X1 U909 ( .A(n1009), .B(n1008), .Y(n1119) );
  NOR3X1 U910 ( .A(sigma3[12]), .B(sigma3[10]), .C(sigma3[11]), .Y(n1008) );
  NOR3X1 U911 ( .A(sigma3[9]), .B(sigma3[7]), .C(sigma3[8]), .Y(n1009) );
  NAND2X1 U912 ( .A(n993), .B(n992), .Y(n997) );
  NOR2X1 U913 ( .A(n1658), .B(sigma15[4]), .Y(n1054) );
  NOR2X1 U914 ( .A(sigma15[11]), .B(sigma15[10]), .Y(n1055) );
  INVX1 U915 ( .A(n1324), .Y(n1370) );
  CLKINVX3 U916 ( .A(n1434), .Y(n1368) );
  OAI21XL U917 ( .A0(n812), .A1(n1386), .B0(n1385), .Y(n1422) );
  NAND2X2 U918 ( .A(n942), .B(n829), .Y(n944) );
  NAND2X1 U919 ( .A(n142), .B(n199), .Y(n235) );
  OAI21X2 U920 ( .A0(n1438), .A1(n881), .B0(n1436), .Y(n1461) );
  AND2X2 U921 ( .A(n214), .B(n815), .Y(n210) );
  AND3X2 U922 ( .A(n1506), .B(n816), .C(n208), .Y(n214) );
  INVX1 U923 ( .A(n1309), .Y(n863) );
  NOR3X1 U924 ( .A(N258), .B(N256), .C(N257), .Y(n1150) );
  CLKINVX3 U925 ( .A(n947), .Y(n948) );
  INVX1 U926 ( .A(n1655), .Y(n1139) );
  NOR3X1 U927 ( .A(sigma6[6]), .B(sigma6[4]), .C(sigma6[5]), .Y(n1071) );
  INVX1 U928 ( .A(n1657), .Y(n852) );
  INVX1 U929 ( .A(n1656), .Y(n854) );
  INVX1 U930 ( .A(n1653), .Y(n845) );
  INVX1 U931 ( .A(n1651), .Y(n848) );
  BUFX3 U932 ( .A(n1650), .Y(sigma11[4]) );
  INVX1 U933 ( .A(n1647), .Y(n834) );
  INVX1 U934 ( .A(n1644), .Y(n843) );
  INVX1 U935 ( .A(N257), .Y(n936) );
  INVXL U936 ( .A(n976), .Y(error_number[0]) );
  INVXL U937 ( .A(n936), .Y(error_number[1]) );
  INVX1 U938 ( .A(n1392), .Y(enable_cs) );
  INVX1 U939 ( .A(n1392), .Y(n1676) );
  NOR2XL U940 ( .A(n1440), .B(n969), .Y(n1442) );
  NOR3X1 U941 ( .A(sigma1[6]), .B(sigma1[4]), .C(n1645), .Y(n1075) );
  INVX1 U942 ( .A(n1649), .Y(n825) );
  INVX1 U943 ( .A(n825), .Y(sigma11[6]) );
  NAND3X1 U944 ( .A(n1065), .B(n1064), .C(n1063), .Y(n1117) );
  NAND2X1 U945 ( .A(n995), .B(n994), .Y(n996) );
  NOR2X1 U946 ( .A(n997), .B(n996), .Y(n1118) );
  INVX1 U947 ( .A(n1321), .Y(n1319) );
  NAND2XL U948 ( .A(n1394), .B(n1384), .Y(n1334) );
  NAND2XL U949 ( .A(sig_all_zero), .B(n1342), .Y(n1407) );
  NAND2XL U950 ( .A(n1340), .B(sig_all_zero), .Y(n1408) );
  AND2X2 U951 ( .A(n1406), .B(n1405), .Y(n828) );
  CLKINVX3 U952 ( .A(n1388), .Y(n1352) );
  XOR3X4 U953 ( .A(n1470), .B(n1471), .C(n1469), .Y(n1457) );
  NAND2XL U954 ( .A(n1431), .B(n1433), .Y(n1355) );
  MX2X4 U955 ( .A(e8), .B(n1312), .S0(n842), .Y(n1363) );
  NOR2X1 U956 ( .A(n1412), .B(n1411), .Y(n829) );
  NOR2X1 U957 ( .A(n1379), .B(n1411), .Y(n1380) );
  NOR3XL U958 ( .A(sigma7[9]), .B(sigma7[7]), .C(sigma7[8]), .Y(n999) );
  INVX2 U959 ( .A(n1413), .Y(n942) );
  NOR3X1 U960 ( .A(sigma9[7]), .B(sigma9[6]), .C(sigma9[8]), .Y(n1062) );
  INVX1 U961 ( .A(n1648), .Y(n830) );
  INVX1 U962 ( .A(n830), .Y(sigma9[3]) );
  NOR3X2 U963 ( .A(sigma10[12]), .B(sigma10[10]), .C(sigma10[11]), .Y(n1000)
         );
  NOR2X2 U964 ( .A(n870), .B(sigma9[11]), .Y(n1061) );
  OAI2BB1XL U965 ( .A0N(n974), .A1N(n1456), .B0(n1455), .Y(n1479) );
  AOI21X1 U966 ( .A0(n1459), .A1(n1468), .B0(n1462), .Y(n1456) );
  BUFX2 U967 ( .A(n1645), .Y(sigma1[5]) );
  NOR3X2 U968 ( .A(sigma2[11]), .B(sigma2[12]), .C(sigma2[10]), .Y(n1032) );
  INVX1 U969 ( .A(n1067), .Y(sigma11[2]) );
  INVX1 U970 ( .A(n834), .Y(sigma9[5]) );
  BUFX2 U971 ( .A(n1646), .Y(sigma2[6]) );
  BUFX2 U972 ( .A(n1323), .Y(n837) );
  INVX1 U973 ( .A(n838), .Y(n839) );
  XNOR2X2 U974 ( .A(n941), .B(n1366), .Y(n1365) );
  NOR3XL U975 ( .A(sigma7[12]), .B(sigma7[10]), .C(sigma7[11]), .Y(n998) );
  NAND2XL U976 ( .A(n1340), .B(sig_all_zero), .Y(n1397) );
  INVX1 U977 ( .A(n1139), .Y(sigma14[11]) );
  NAND4XL U978 ( .A(n1013), .B(n1012), .C(n1011), .D(n1010), .Y(n841) );
  NOR2X2 U979 ( .A(sigma2[6]), .B(sigma2[4]), .Y(n1011) );
  NAND2X2 U980 ( .A(n1507), .B(n1340), .Y(n874) );
  CLKINVX3 U981 ( .A(n884), .Y(n941) );
  NAND2X2 U982 ( .A(n876), .B(n877), .Y(n879) );
  NAND2X2 U983 ( .A(n878), .B(n879), .Y(n1361) );
  INVX1 U984 ( .A(n1652), .Y(n1067) );
  MXI2X1 U985 ( .A(n900), .B(n1305), .S0(n1345), .Y(n884) );
  INVX1 U986 ( .A(sigma11[7]), .Y(n1064) );
  XOR2X2 U987 ( .A(n1354), .B(n1353), .Y(n1429) );
  NOR2X1 U988 ( .A(sigma14[2]), .B(n1656), .Y(n1057) );
  AND2X4 U989 ( .A(n1376), .B(n1375), .Y(n873) );
  NAND2X1 U990 ( .A(n602), .B(n875), .Y(n1403) );
  INVX1 U991 ( .A(n843), .Y(sigma1[8]) );
  INVX1 U992 ( .A(n845), .Y(sigma11[1]) );
  BUFX2 U993 ( .A(n1654), .Y(sigma12[4]) );
  OAI21X1 U994 ( .A0(n1395), .A1(n1506), .B0(n1394), .Y(n1399) );
  NAND2X2 U995 ( .A(n1482), .B(n1490), .Y(n1441) );
  INVX1 U996 ( .A(n848), .Y(sigma11[3]) );
  MXI2X1 U997 ( .A(n594), .B(n1115), .S0(n1345), .Y(n1362) );
  XNOR2X2 U998 ( .A(n1457), .B(n1458), .Y(n1500) );
  MXI2X4 U999 ( .A(n597), .B(n1134), .S0(n1345), .Y(n1411) );
  OR2X4 U1000 ( .A(n1431), .B(n1429), .Y(n1460) );
  NAND2X2 U1001 ( .A(n1374), .B(n1375), .Y(n1382) );
  OAI22X1 U1002 ( .A0(n941), .A1(n839), .B0(n1365), .B1(n1364), .Y(n1434) );
  NAND2X1 U1003 ( .A(n1404), .B(n1403), .Y(n1389) );
  NAND2X2 U1004 ( .A(n1345), .B(n1344), .Y(n1404) );
  NOR4X2 U1005 ( .A(sigma10[2]), .B(sigma10[3]), .C(sigma10[0]), .D(sigma10[1]), .Y(n1003) );
  OR2X2 U1006 ( .A(err_count[8]), .B(err_count[7]), .Y(n980) );
  NAND4X2 U1007 ( .A(n850), .B(n1035), .C(n1037), .D(n1036), .Y(n1038) );
  NAND2X4 U1008 ( .A(n1329), .B(n1328), .Y(sig_all_zero) );
  NOR2X1 U1009 ( .A(sigma11[9]), .B(sigma11[12]), .Y(n1063) );
  CLKINVX3 U1010 ( .A(n1327), .Y(n1081) );
  NAND4X2 U1011 ( .A(n1080), .B(n1079), .C(n1078), .D(n1077), .Y(n1327) );
  NOR4BX2 U1012 ( .AN(n1034), .B(n1123), .C(n1122), .D(n1125), .Y(n1035) );
  CLKINVX4 U1013 ( .A(n1038), .Y(n1329) );
  NOR3X2 U1014 ( .A(sigma1[9]), .B(sigma1[7]), .C(n1644), .Y(n1074) );
  NOR2X1 U1015 ( .A(err_count[11]), .B(err_count[9]), .Y(n978) );
  NOR3X2 U1016 ( .A(n1305), .B(n1120), .C(n1119), .Y(n1037) );
  CLKINVX8 U1017 ( .A(n1103), .Y(n1328) );
  INVX1 U1018 ( .A(n852), .Y(sigma14[0]) );
  INVX1 U1019 ( .A(n854), .Y(sigma14[1]) );
  INVX2 U1020 ( .A(n1379), .Y(n1375) );
  NAND2X1 U1021 ( .A(n1318), .B(n1317), .Y(n1321) );
  NAND2X1 U1022 ( .A(n817), .B(n1345), .Y(n1318) );
  INVX1 U1023 ( .A(n856), .Y(n857) );
  INVX1 U1024 ( .A(n890), .Y(n858) );
  INVX1 U1025 ( .A(n893), .Y(n859) );
  INVX1 U1026 ( .A(n895), .Y(n860) );
  INVX1 U1027 ( .A(n1675), .Y(n861) );
  INVX1 U1028 ( .A(n861), .Y(count[5]) );
  INVX1 U1029 ( .A(n894), .Y(n864) );
  OAI22XL U1030 ( .A0(n580), .A1(n124), .B0(n86), .B1(n125), .Y(n704) );
  OAI22XL U1031 ( .A0(n581), .A1(n124), .B0(n87), .B1(n125), .Y(n705) );
  INVX1 U1032 ( .A(n891), .Y(n865) );
  OAI22XL U1033 ( .A0(n555), .A1(n116), .B0(n87), .B1(n117), .Y(n679) );
  OAI22XL U1034 ( .A0(n554), .A1(n116), .B0(n86), .B1(n117), .Y(n678) );
  INVX1 U1035 ( .A(n892), .Y(n866) );
  OAI22XL U1036 ( .A0(n530), .A1(n107), .B0(n87), .B1(n108), .Y(n654) );
  OAI22XL U1037 ( .A0(n531), .A1(n107), .B0(n86), .B1(n108), .Y(n655) );
  INVX1 U1038 ( .A(n888), .Y(n867) );
  OAI22XL U1039 ( .A0(n489), .A1(n79), .B0(n86), .B1(n81), .Y(n613) );
  OAI22XL U1040 ( .A0(n490), .A1(n79), .B0(n87), .B1(n81), .Y(n614) );
  OAI22XL U1041 ( .A0(n518), .A1(n1504), .B0(n86), .B1(n949), .Y(n642) );
  OAI22XL U1042 ( .A0(n517), .A1(n1504), .B0(n87), .B1(n949), .Y(n641) );
  INVX1 U1043 ( .A(n896), .Y(n868) );
  NAND2XL U1044 ( .A(N670), .B(n868), .Y(n131) );
  AOI22XL U1045 ( .A0(err_count[12]), .A1(n127), .B0(N661), .B1(n128), .Y(n85)
         );
  AOI22XL U1046 ( .A0(n951), .A1(err_count[11]), .B0(N662), .B1(n128), .Y(n90)
         );
  AOI22XL U1047 ( .A0(n951), .A1(err_count[7]), .B0(N666), .B1(n128), .Y(n88)
         );
  NOR3X1 U1048 ( .A(n970), .B(n868), .C(n195), .Y(n196) );
  NOR3X2 U1049 ( .A(sigma1[12]), .B(sigma1[10]), .C(sigma1[11]), .Y(n1073) );
  NOR2X1 U1050 ( .A(sigma16[0]), .B(sigma16[11]), .Y(n1051) );
  OAI21X1 U1051 ( .A0(n1393), .A1(n1392), .B0(n763), .Y(n1405) );
  NAND2X1 U1052 ( .A(n1107), .B(n1106), .Y(n871) );
  NOR2XL U1053 ( .A(sigma15[4]), .B(sigma15[3]), .Y(n1110) );
  NAND2X2 U1054 ( .A(n1106), .B(n1107), .Y(n1338) );
  NAND2XL U1055 ( .A(n1394), .B(n1384), .Y(n1385) );
  NAND2BX1 U1056 ( .AN(n1367), .B(n882), .Y(n1437) );
  NOR2X2 U1057 ( .A(n819), .B(n1130), .Y(n1100) );
  XNOR3X4 U1058 ( .A(n1382), .B(n873), .C(n1381), .Y(n1458) );
  NOR4X2 U1059 ( .A(sigma6[2]), .B(sigma6[3]), .C(sigma6[0]), .D(sigma6[1]), 
        .Y(n1072) );
  NOR2X2 U1060 ( .A(n818), .B(n1058), .Y(n1101) );
  NAND3X2 U1061 ( .A(n1102), .B(n1100), .C(n1101), .Y(n947) );
  NOR2XL U1062 ( .A(n1657), .B(sigma15[12]), .Y(n1056) );
  OAI2BB1XL U1063 ( .A0N(n1493), .A1N(n1492), .B0(n1491), .Y(n1499) );
  INVX1 U1064 ( .A(n1362), .Y(n876) );
  NOR2X1 U1065 ( .A(n1150), .B(n1277), .Y(n977) );
  NOR4X2 U1066 ( .A(sigma1[2]), .B(sigma1[3]), .C(sigma1[0]), .D(sigma1[1]), 
        .Y(n1076) );
  INVXL U1067 ( .A(n1437), .Y(n880) );
  XNOR2X1 U1068 ( .A(n1361), .B(n1313), .Y(n882) );
  NAND2XL U1069 ( .A(n1362), .B(n1363), .Y(n878) );
  INVX1 U1070 ( .A(n1363), .Y(n877) );
  OAI22X1 U1071 ( .A0(n1363), .A1(n1362), .B0(n1361), .B1(n1360), .Y(n1435) );
  OAI21X1 U1072 ( .A0(n1471), .A1(n1453), .B0(n1452), .Y(n1443) );
  OR2XL U1073 ( .A(n1132), .B(n1133), .Y(n1295) );
  NOR2X1 U1074 ( .A(sigma13[4]), .B(sigma13[5]), .Y(n1086) );
  NAND2X1 U1075 ( .A(n1422), .B(n1421), .Y(n1453) );
  NOR2X1 U1076 ( .A(n980), .B(n981), .Y(n898) );
  NAND2X2 U1077 ( .A(n1096), .B(n1095), .Y(n1097) );
  NAND3X1 U1078 ( .A(n1503), .B(n1502), .C(n1501), .Y(n1508) );
  NAND2BX1 U1079 ( .AN(err_count[5]), .B(n898), .Y(n983) );
  INVXL U1080 ( .A(sigma14[4]), .Y(n1039) );
  NAND3BXL U1081 ( .AN(sigma14[2]), .B(n1136), .C(n1135), .Y(n1288) );
  NOR2XL U1082 ( .A(sigma14[3]), .B(sigma14[4]), .Y(n1136) );
  NOR2XL U1083 ( .A(sigma15[1]), .B(sigma15[0]), .Y(n1109) );
  NAND3XL U1084 ( .A(n1355), .B(n1460), .C(n1416), .Y(n1427) );
  NAND2BXL U1085 ( .AN(n1494), .B(n1490), .Y(n1481) );
  NOR3XL U1086 ( .A(n1485), .B(n1484), .C(n1493), .Y(n1486) );
  NAND2XL U1087 ( .A(n967), .B(n811), .Y(n1495) );
  INVXL U1088 ( .A(n1482), .Y(n1480) );
  NAND2BX1 U1089 ( .AN(n1500), .B(n1491), .Y(n1440) );
  INVXL U1090 ( .A(n1460), .Y(n1472) );
  NAND3BXL U1091 ( .AN(n1433), .B(n1432), .C(n1473), .Y(n1490) );
  INVXL U1092 ( .A(n1431), .Y(n1432) );
  AOI21XL U1093 ( .A0(n1472), .A1(n1473), .B0(n1461), .Y(n1464) );
  INVXL U1094 ( .A(n1461), .Y(n1493) );
  OAI2BB1X1 U1095 ( .A0N(n886), .A1N(n1469), .B0(n1454), .Y(n1462) );
  INVX1 U1096 ( .A(n1357), .Y(n1416) );
  NOR2XL U1097 ( .A(n1341), .B(n871), .Y(n1342) );
  NAND2XL U1098 ( .A(n1422), .B(n1421), .Y(n1470) );
  NAND2BXL U1099 ( .AN(n1473), .B(n1380), .Y(n946) );
  INVX2 U1100 ( .A(n1435), .Y(n1369) );
  NOR2X4 U1101 ( .A(n1098), .B(n1097), .Y(n1099) );
  XOR2X1 U1102 ( .A(n1367), .B(n882), .Y(n1357) );
  INVX1 U1103 ( .A(n1308), .Y(n1315) );
  AOI211X1 U1104 ( .A0(N672), .A1(n128), .B0(n137), .C0(n138), .Y(n136) );
  NAND2X1 U1105 ( .A(n967), .B(n144), .Y(n92) );
  NAND2XL U1106 ( .A(n1121), .B(n883), .Y(n1332) );
  NAND2XL U1107 ( .A(n1118), .B(n885), .Y(n1311) );
  INVXL U1108 ( .A(n1320), .Y(n1322) );
  NOR2X1 U1109 ( .A(n206), .B(n821), .Y(n212) );
  XNOR2X1 U1110 ( .A(n1365), .B(n1364), .Y(n1367) );
  OR2XL U1111 ( .A(n1143), .B(n1144), .Y(n1291) );
  OR2XL U1112 ( .A(n1117), .B(n1116), .Y(n1301) );
  OR2XL U1113 ( .A(n1104), .B(n1105), .Y(n1151) );
  NOR2XL U1114 ( .A(n1131), .B(n1308), .Y(n1147) );
  NAND3XL U1115 ( .A(n1147), .B(n1411), .C(n1146), .Y(n1148) );
  AOI22XL U1116 ( .A0(n951), .A1(err_count[10]), .B0(N663), .B1(n128), .Y(n86)
         );
  AOI22XL U1117 ( .A0(n951), .A1(err_count[8]), .B0(N665), .B1(n128), .Y(n87)
         );
  NOR3XL U1118 ( .A(sigma13[11]), .B(n1291), .C(n1292), .Y(n1145) );
  AND2X2 U1119 ( .A(n991), .B(n990), .Y(n883) );
  OAI2BB1X1 U1120 ( .A0N(n130), .A1N(n131), .B0(n973), .Y(n83) );
  NAND3X1 U1121 ( .A(n1016), .B(n1015), .C(n1014), .Y(n1133) );
  INVXL U1122 ( .A(sigma12[2]), .Y(n1015) );
  NAND3X1 U1123 ( .A(n1094), .B(n1093), .C(n1092), .Y(n1104) );
  INVXL U1124 ( .A(sigma16[2]), .Y(n1093) );
  NAND3X1 U1125 ( .A(n1088), .B(n1087), .C(n1086), .Y(n1143) );
  NOR2XL U1126 ( .A(sigma14[3]), .B(sigma14[5]), .Y(n1040) );
  NAND2XL U1127 ( .A(n1355), .B(n1460), .Y(n1356) );
  NAND4X1 U1128 ( .A(n1029), .B(n1028), .C(n1027), .D(n1026), .Y(n1123) );
  NAND4X1 U1129 ( .A(n1007), .B(n1006), .C(n1005), .D(n1004), .Y(n1120) );
  NAND3X1 U1130 ( .A(n1019), .B(n1018), .C(n1017), .Y(n1132) );
  NOR2XL U1131 ( .A(n1655), .B(sigma14[10]), .Y(n1041) );
  NAND3BXL U1132 ( .AN(sigma15[2]), .B(n1110), .C(n1109), .Y(n1281) );
  NOR2X1 U1133 ( .A(sigma8[4]), .B(sigma8[5]), .Y(n1026) );
  NOR2X1 U1134 ( .A(sigma3[4]), .B(sigma3[5]), .Y(n1004) );
  NAND3X1 U1135 ( .A(n1091), .B(n1090), .C(n1089), .Y(n1105) );
  INVXL U1136 ( .A(sigma16[7]), .Y(n1090) );
  NAND3X1 U1137 ( .A(n1085), .B(n1084), .C(n1083), .Y(n1144) );
  INVXL U1138 ( .A(sigma13[7]), .Y(n1084) );
  NOR2XL U1139 ( .A(sigma14[7]), .B(sigma14[6]), .Y(n1138) );
  NOR2XL U1140 ( .A(sigma14[9]), .B(sigma14[8]), .Y(n1137) );
  NOR2XL U1141 ( .A(sigma15[7]), .B(sigma15[6]), .Y(n1112) );
  NOR2XL U1142 ( .A(sigma15[9]), .B(sigma15[8]), .Y(n1111) );
  INVXL U1143 ( .A(sigma14[12]), .Y(n1286) );
  NAND2XL U1144 ( .A(n1487), .B(n1476), .Y(n1477) );
  NAND2X1 U1145 ( .A(n1031), .B(n1030), .Y(n1122) );
  AOI221XL U1146 ( .A0(n110), .A1(n157), .B0(n155), .B1(N257), .C0(n114), .Y(
        n156) );
  OR2XL U1147 ( .A(sigma13[10]), .B(sigma13[0]), .Y(n1292) );
  OR2XL U1148 ( .A(sigma12[10]), .B(sigma12[0]), .Y(n1296) );
  NAND2X1 U1149 ( .A(n1046), .B(n1045), .Y(n1047) );
  NOR2XL U1150 ( .A(sigma11[11]), .B(sigma11[10]), .Y(n1046) );
  NOR2XL U1151 ( .A(sigma11[0]), .B(sigma12[11]), .Y(n1045) );
  OR2XL U1152 ( .A(sigma16[0]), .B(sigma16[10]), .Y(n1152) );
  OR2XL U1153 ( .A(sigma15[10]), .B(sigma15[5]), .Y(n1113) );
  OR2XL U1154 ( .A(sigma14[10]), .B(sigma14[5]), .Y(n1140) );
  AND2X2 U1155 ( .A(n999), .B(n998), .Y(n885) );
  NOR2XL U1156 ( .A(n976), .B(N257), .Y(n110) );
  AOI21XL U1157 ( .A0(n142), .A1(n874), .B0(n1315), .Y(n1310) );
  NOR2XL U1158 ( .A(n936), .B(N256), .Y(n114) );
  NOR2XL U1159 ( .A(n195), .B(error_number[3]), .Y(n106) );
  INVXL U1160 ( .A(N256), .Y(n976) );
  NOR2XL U1161 ( .A(n1296), .B(sigma12[11]), .Y(n1297) );
  INVXL U1162 ( .A(N258), .Y(n115) );
  AND2X1 U1163 ( .A(n106), .B(N258), .Y(n101) );
  NOR4BXL U1164 ( .AN(n856), .B(n1292), .C(sigma13[11]), .D(n1291), .Y(n1293)
         );
  NOR4BXL U1165 ( .AN(n856), .B(n1302), .C(sigma11[11]), .D(n1301), .Y(n1303)
         );
  NOR3XL U1166 ( .A(sigma14[5]), .B(n1655), .C(sigma14[10]), .Y(n1285) );
  NOR3XL U1167 ( .A(sigma15[5]), .B(sigma15[11]), .C(sigma15[10]), .Y(n1278)
         );
  NAND2XL U1168 ( .A(n970), .B(e_sum_r[2]), .Y(n1445) );
  CLKBUFXL U1169 ( .A(error_number[3]), .Y(serr[3]) );
  CLKBUFXL U1170 ( .A(N258), .Y(error_number[2]) );
  INVX1 U1171 ( .A(n1494), .Y(n1483) );
  INVX1 U1172 ( .A(n965), .Y(n963) );
  INVX1 U1173 ( .A(n965), .Y(n962) );
  INVX1 U1174 ( .A(n966), .Y(n961) );
  INVX1 U1175 ( .A(n966), .Y(n960) );
  INVX1 U1176 ( .A(n966), .Y(n959) );
  INVX1 U1177 ( .A(n966), .Y(n957) );
  INVX1 U1178 ( .A(n966), .Y(n956) );
  INVX1 U1179 ( .A(n966), .Y(n955) );
  INVX1 U1180 ( .A(n966), .Y(n958) );
  INVX1 U1181 ( .A(n966), .Y(n953) );
  INVX1 U1182 ( .A(n966), .Y(n954) );
  INVX1 U1183 ( .A(n965), .Y(n964) );
  INVX1 U1184 ( .A(n1309), .Y(n1300) );
  NAND2X1 U1185 ( .A(n967), .B(n1483), .Y(n1488) );
  NAND2X1 U1186 ( .A(n967), .B(n1444), .Y(n1455) );
  NOR2X1 U1187 ( .A(n1481), .B(n1480), .Y(n1485) );
  NAND3X1 U1188 ( .A(n1467), .B(n1466), .C(n1491), .Y(n1478) );
  NAND3X1 U1189 ( .A(n1465), .B(n1464), .C(n1463), .Y(n1466) );
  INVXL U1190 ( .A(n1462), .Y(n1463) );
  INVX1 U1191 ( .A(n887), .Y(n965) );
  INVX1 U1192 ( .A(n79), .Y(n81) );
  INVX1 U1193 ( .A(n887), .Y(n966) );
  OAI21XL U1194 ( .A0(n1474), .A1(n1473), .B0(n1472), .Y(n1497) );
  INVX1 U1195 ( .A(n1489), .Y(n1474) );
  XOR3X2 U1196 ( .A(n1369), .B(n1368), .C(n881), .Y(n1426) );
  OAI21XL U1197 ( .A0(n1429), .A1(n1431), .B0(n1428), .Y(n1459) );
  OR2X2 U1198 ( .A(n1471), .B(n1470), .Y(n886) );
  NAND2X2 U1199 ( .A(n1430), .B(n1459), .Y(n1482) );
  XOR3X2 U1200 ( .A(n1453), .B(n1471), .C(n1452), .Y(n1430) );
  NAND2X1 U1201 ( .A(n945), .B(n946), .Y(n1381) );
  XNOR3X2 U1202 ( .A(n1369), .B(n1368), .C(n1437), .Y(n940) );
  XOR3X2 U1203 ( .A(n1494), .B(n1461), .C(n1441), .Y(n1439) );
  NAND3X1 U1204 ( .A(n1417), .B(n1460), .C(n1416), .Y(n1418) );
  AND2X2 U1205 ( .A(n967), .B(n1676), .Y(n887) );
  INVX1 U1206 ( .A(n971), .Y(n967) );
  XOR2X1 U1207 ( .A(n1453), .B(n1471), .Y(n1419) );
  OR2X2 U1208 ( .A(n970), .B(n82), .Y(n888) );
  INVX1 U1209 ( .A(n888), .Y(n79) );
  INVX1 U1210 ( .A(n116), .Y(n117) );
  INVX1 U1211 ( .A(n121), .Y(n122) );
  INVX1 U1212 ( .A(n98), .Y(n99) );
  INVX1 U1213 ( .A(n107), .Y(n108) );
  INVX1 U1214 ( .A(n111), .Y(n112) );
  INVX1 U1215 ( .A(n124), .Y(n125) );
  INVX1 U1216 ( .A(n949), .Y(n1504) );
  INVX1 U1217 ( .A(n971), .Y(n968) );
  NOR3X1 U1218 ( .A(n211), .B(n145), .C(n212), .Y(n198) );
  NAND2X1 U1219 ( .A(n1415), .B(n1414), .Y(n1424) );
  NAND3X1 U1220 ( .A(n1371), .B(n1378), .C(n1370), .Y(n1377) );
  INVX1 U1221 ( .A(n1389), .Y(n1350) );
  XNOR3X2 U1222 ( .A(n1352), .B(n889), .C(n1389), .Y(n1415) );
  NAND3X1 U1223 ( .A(n1371), .B(n1378), .C(n1370), .Y(n1372) );
  XOR3X2 U1224 ( .A(n1352), .B(n1351), .C(n1350), .Y(n1353) );
  XNOR3X2 U1225 ( .A(n1402), .B(n812), .C(n1349), .Y(n1354) );
  NAND3X1 U1226 ( .A(n1451), .B(n1450), .C(n1449), .Y(n1509) );
  NAND3X1 U1227 ( .A(n1448), .B(n1447), .C(n1446), .Y(n1449) );
  INVX1 U1228 ( .A(n196), .Y(n155) );
  INVX1 U1229 ( .A(n1343), .Y(n1344) );
  INVX1 U1230 ( .A(n1321), .Y(n1314) );
  INVX1 U1231 ( .A(n972), .Y(n971) );
  NAND2X1 U1232 ( .A(n96), .B(n97), .Y(n82) );
  OR2X2 U1233 ( .A(n970), .B(n123), .Y(n890) );
  INVX1 U1234 ( .A(n890), .Y(n121) );
  OR2X2 U1235 ( .A(n970), .B(n118), .Y(n891) );
  INVX1 U1236 ( .A(n891), .Y(n116) );
  INVX1 U1237 ( .A(n97), .Y(n153) );
  OR2X2 U1238 ( .A(n969), .B(n109), .Y(n892) );
  INVX1 U1239 ( .A(n892), .Y(n107) );
  OR2X2 U1240 ( .A(n970), .B(n113), .Y(n893) );
  INVX1 U1241 ( .A(n893), .Y(n111) );
  OR2X2 U1242 ( .A(n970), .B(n129), .Y(n894) );
  INVX1 U1243 ( .A(n894), .Y(n124) );
  OR2X2 U1244 ( .A(n970), .B(n100), .Y(n895) );
  INVX1 U1245 ( .A(n895), .Y(n98) );
  INVX1 U1246 ( .A(n973), .Y(n970) );
  BUFX3 U1247 ( .A(n1629), .Y(n949) );
  NAND2BX1 U1248 ( .AN(n1156), .B(n967), .Y(n1629) );
  INVX1 U1249 ( .A(n974), .Y(n969) );
  NAND2X1 U1250 ( .A(n1312), .B(n1343), .Y(n1126) );
  INVX1 U1251 ( .A(n72), .Y(pre_err) );
  NOR2X1 U1252 ( .A(n1025), .B(n1024), .Y(n1034) );
  NAND2X1 U1253 ( .A(n1021), .B(n1020), .Y(n1025) );
  NAND2X1 U1254 ( .A(n1023), .B(n1022), .Y(n1024) );
  MX2X1 U1255 ( .A(n910), .B(n909), .S0(error_number[2]), .Y(N672) );
  NAND4X1 U1256 ( .A(n198), .B(n165), .C(n175), .D(n135), .Y(n143) );
  OAI21XL U1257 ( .A0(n1389), .A1(n1390), .B0(n1388), .Y(n1423) );
  NAND3X1 U1258 ( .A(n814), .B(n822), .C(n225), .Y(n206) );
  NOR2X1 U1259 ( .A(n235), .B(n820), .Y(n145) );
  AOI21X2 U1260 ( .A0(n837), .A1(n1320), .B0(n1314), .Y(n1326) );
  NOR3BX2 U1261 ( .AN(n1323), .B(n1316), .C(n1322), .Y(n1325) );
  OR2XL U1262 ( .A(n841), .B(n1125), .Y(n1343) );
  NAND3X1 U1263 ( .A(n133), .B(n146), .C(n77), .Y(n197) );
  NAND2X1 U1264 ( .A(n1406), .B(n1405), .Y(n1388) );
  NAND2X1 U1265 ( .A(n1323), .B(n1320), .Y(n1308) );
  INVX1 U1266 ( .A(n1360), .Y(n1313) );
  XOR2X1 U1267 ( .A(n1348), .B(n1347), .Y(n1349) );
  NAND4BXL U1268 ( .AN(n145), .B(n146), .C(n147), .D(n148), .Y(n144) );
  AOI211X1 U1269 ( .A0(N671), .A1(n128), .B0(n137), .C0(n149), .Y(n148) );
  MX2X1 U1270 ( .A(n912), .B(n911), .S0(error_number[2]), .Y(N671) );
  INVX1 U1271 ( .A(n147), .Y(n172) );
  XOR3X2 U1272 ( .A(n1400), .B(n1335), .C(n1334), .Y(n1414) );
  NAND2X1 U1273 ( .A(n1383), .B(n1396), .Y(n1335) );
  INVX1 U1274 ( .A(n134), .Y(n211) );
  OR2XL U1275 ( .A(n1119), .B(n1120), .Y(n1341) );
  OAI21XL U1276 ( .A0(n1277), .A1(n192), .B0(n194), .Y(n736) );
  NOR3X1 U1277 ( .A(n155), .B(n153), .C(n115), .Y(n192) );
  OR4X2 U1278 ( .A(n897), .B(n143), .C(n197), .D(n137), .Y(n896) );
  OR3XL U1279 ( .A(n138), .B(n172), .C(n160), .Y(n897) );
  OAI2BB1X1 U1280 ( .A0N(n1488), .A1N(n1487), .B0(n1486), .Y(n1502) );
  OAI211X1 U1281 ( .A0(n199), .A1(n204), .B0(n813), .C0(n823), .Y(n137) );
  INVX1 U1282 ( .A(n976), .Y(n935) );
  INVX1 U1283 ( .A(n976), .Y(n934) );
  NOR2X1 U1284 ( .A(n1144), .B(n1143), .Y(n1096) );
  INVX1 U1285 ( .A(n200), .Y(n160) );
  BUFX3 U1286 ( .A(n127), .Y(n951) );
  NAND4BXL U1287 ( .AN(n197), .B(n198), .C(n130), .D(n199), .Y(n127) );
  INVX1 U1288 ( .A(n182), .Y(n1505) );
  OR2XL U1289 ( .A(n1122), .B(n1123), .Y(n1312) );
  INVX1 U1290 ( .A(n975), .Y(n972) );
  NOR4BX1 U1291 ( .AN(n256), .B(count[5]), .C(count[6]), .D(n952), .Y(n253) );
  NAND3X1 U1292 ( .A(n976), .B(n936), .C(n101), .Y(n118) );
  NOR2X1 U1293 ( .A(n936), .B(n976), .Y(n97) );
  AOI21X1 U1294 ( .A0(n133), .A1(n874), .B0(n971), .Y(n1284) );
  NAND2X1 U1295 ( .A(n110), .B(n101), .Y(n123) );
  NAND2X1 U1296 ( .A(n101), .B(n97), .Y(n100) );
  NAND2X1 U1297 ( .A(n110), .B(n96), .Y(n109) );
  NAND2X1 U1298 ( .A(n114), .B(n96), .Y(n113) );
  NAND2X1 U1299 ( .A(n114), .B(n101), .Y(n129) );
  NAND2X1 U1300 ( .A(N264), .B(N263), .Y(n251) );
  NAND4BXL U1301 ( .AN(count[2]), .B(n253), .C(n254), .D(n255), .Y(n248) );
  MXI2X1 U1302 ( .A(n1269), .B(n1270), .S0(n953), .Y(n1516) );
  MXI2X1 U1303 ( .A(n1195), .B(n1196), .S0(n960), .Y(n1591) );
  MXI2X1 U1304 ( .A(n1172), .B(n1173), .S0(n962), .Y(n1614) );
  MXI2X1 U1305 ( .A(n1196), .B(n1197), .S0(n960), .Y(n1590) );
  MXI2X1 U1306 ( .A(n1262), .B(n1264), .S0(n953), .Y(n1523) );
  MXI2X1 U1307 ( .A(n1266), .B(n1267), .S0(n953), .Y(n1519) );
  MXI2X1 U1308 ( .A(n1234), .B(n1235), .S0(n956), .Y(n1551) );
  MXI2X1 U1309 ( .A(n1205), .B(n1206), .S0(n959), .Y(n1581) );
  MXI2X1 U1310 ( .A(n1179), .B(n1180), .S0(n961), .Y(n1607) );
  MXI2X1 U1311 ( .A(n1214), .B(n1215), .S0(n958), .Y(n1572) );
  MXI2X1 U1312 ( .A(n1217), .B(n1218), .S0(n958), .Y(n1569) );
  MXI2X1 U1313 ( .A(n1241), .B(n1242), .S0(n955), .Y(n1544) );
  MXI2X1 U1314 ( .A(n1243), .B(n1244), .S0(n955), .Y(n1542) );
  MXI2X1 U1315 ( .A(n1165), .B(n1166), .S0(n962), .Y(n1625) );
  MXI2X1 U1316 ( .A(n1169), .B(n1170), .S0(n962), .Y(n1617) );
  MXI2X1 U1317 ( .A(n1170), .B(n1171), .S0(n961), .Y(n1616) );
  MXI2X1 U1318 ( .A(n1178), .B(n1179), .S0(n961), .Y(n1608) );
  MXI2X1 U1319 ( .A(n1181), .B(n1182), .S0(n961), .Y(n1605) );
  MXI2X1 U1320 ( .A(n1182), .B(n1184), .S0(n961), .Y(n1604) );
  MXI2X1 U1321 ( .A(n1186), .B(n1187), .S0(n961), .Y(n1600) );
  MXI2X1 U1322 ( .A(n1197), .B(n1198), .S0(n959), .Y(n1589) );
  MXI2X1 U1323 ( .A(n1200), .B(n1202), .S0(n959), .Y(n1586) );
  MXI2X1 U1324 ( .A(n1206), .B(n1207), .S0(n959), .Y(n1580) );
  MXI2X1 U1325 ( .A(n1225), .B(n1226), .S0(n957), .Y(n1560) );
  MXI2X1 U1326 ( .A(n1226), .B(n1228), .S0(n957), .Y(n1559) );
  MXI2X1 U1327 ( .A(n1232), .B(n1233), .S0(n956), .Y(n1553) );
  MXI2X1 U1328 ( .A(n1235), .B(n1237), .S0(n956), .Y(n1550) );
  MXI2X1 U1329 ( .A(n1257), .B(n1258), .S0(n954), .Y(n1528) );
  MXI2X1 U1330 ( .A(n1261), .B(n1262), .S0(n954), .Y(n1524) );
  MXI2X1 U1331 ( .A(n1187), .B(n1188), .S0(n960), .Y(n1599) );
  MXI2X1 U1332 ( .A(n1188), .B(n1189), .S0(n960), .Y(n1598) );
  MXI2X1 U1333 ( .A(n1222), .B(n1223), .S0(n957), .Y(n1563) );
  MXI2X1 U1334 ( .A(n1230), .B(n1231), .S0(n956), .Y(n1555) );
  MXI2X1 U1335 ( .A(n1250), .B(n1251), .S0(n955), .Y(n1535) );
  MXI2X1 U1336 ( .A(n1252), .B(n1253), .S0(n954), .Y(n1533) );
  MXI2X1 U1337 ( .A(n1240), .B(n1241), .S0(n955), .Y(n1545) );
  MXI2X1 U1338 ( .A(n1268), .B(n1269), .S0(n953), .Y(n1517) );
  MXI2X1 U1339 ( .A(n1167), .B(n1168), .S0(n963), .Y(n1623) );
  MXI2X1 U1340 ( .A(n1208), .B(n1209), .S0(n958), .Y(n1578) );
  MXI2X1 U1341 ( .A(n1213), .B(n1214), .S0(n958), .Y(n1573) );
  MXI2X1 U1342 ( .A(n1244), .B(n1246), .S0(n955), .Y(n1541) );
  MXI2X1 U1343 ( .A(n1218), .B(n1220), .S0(n957), .Y(n1568) );
  MXI2X1 U1344 ( .A(n1253), .B(n1255), .S0(n954), .Y(n1532) );
  MXI2X1 U1345 ( .A(n1259), .B(n1260), .S0(n954), .Y(n1526) );
  MXI2X1 U1346 ( .A(n1164), .B(n1165), .S0(n963), .Y(n1626) );
  MXI2X1 U1347 ( .A(n1189), .B(n1190), .S0(n960), .Y(n1597) );
  MXI2X1 U1348 ( .A(n1258), .B(n1259), .S0(n954), .Y(n1527) );
  MXI2X1 U1349 ( .A(n1166), .B(n1167), .S0(n962), .Y(n1624) );
  MXI2X1 U1350 ( .A(n1171), .B(n1172), .S0(n962), .Y(n1615) );
  MXI2X1 U1351 ( .A(n1191), .B(n1193), .S0(n960), .Y(n1595) );
  MXI2X1 U1352 ( .A(n1198), .B(n1199), .S0(n959), .Y(n1588) );
  MXI2X1 U1353 ( .A(n1207), .B(n1208), .S0(n959), .Y(n1579) );
  MXI2X1 U1354 ( .A(n1215), .B(n1216), .S0(n958), .Y(n1571) );
  MXI2X1 U1355 ( .A(n1216), .B(n1217), .S0(n958), .Y(n1570) );
  MXI2X1 U1356 ( .A(n1221), .B(n1222), .S0(n957), .Y(n1564) );
  MXI2X1 U1357 ( .A(n1223), .B(n1224), .S0(n957), .Y(n1562) );
  MXI2X1 U1358 ( .A(n1231), .B(n1232), .S0(n956), .Y(n1554) );
  MXI2X1 U1359 ( .A(n1233), .B(n1234), .S0(n956), .Y(n1552) );
  MXI2X1 U1360 ( .A(n1260), .B(n1261), .S0(n958), .Y(n1525) );
  MXI2X1 U1361 ( .A(n1224), .B(n1225), .S0(n957), .Y(n1561) );
  MXI2X1 U1362 ( .A(n1239), .B(n1240), .S0(n956), .Y(n1546) );
  MXI2X1 U1363 ( .A(n1173), .B(n1175), .S0(n962), .Y(n1613) );
  MXI2X1 U1364 ( .A(n1177), .B(n1178), .S0(n962), .Y(n1609) );
  MXI2X1 U1365 ( .A(n1190), .B(n1191), .S0(n960), .Y(n1596) );
  MXI2X1 U1366 ( .A(n1199), .B(n1200), .S0(n959), .Y(n1587) );
  MXI2X1 U1367 ( .A(n1209), .B(n1211), .S0(n958), .Y(n1577) );
  MXI2X1 U1368 ( .A(n1249), .B(n1250), .S0(n955), .Y(n1536) );
  MXI2X1 U1369 ( .A(n1251), .B(n1252), .S0(n954), .Y(n1534) );
  MXI2X1 U1370 ( .A(n1270), .B(n1271), .S0(n953), .Y(n1515) );
  MXI2X1 U1371 ( .A(n1271), .B(n1273), .S0(n953), .Y(n1514) );
  MXI2X1 U1372 ( .A(n1180), .B(n1181), .S0(n961), .Y(n1606) );
  MXI2X1 U1373 ( .A(n1204), .B(n1205), .S0(n959), .Y(n1582) );
  MXI2X1 U1374 ( .A(n1248), .B(n1249), .S0(n955), .Y(n1537) );
  MXI2X1 U1375 ( .A(n1267), .B(n1268), .S0(n953), .Y(n1518) );
  MXI2X1 U1376 ( .A(n1242), .B(n1243), .S0(n955), .Y(n1543) );
  AND2X2 U1377 ( .A(n106), .B(n115), .Y(n96) );
  AND4X2 U1378 ( .A(count[3]), .B(count[2]), .C(count[1]), .D(n253), .Y(n250)
         );
  INVX1 U1379 ( .A(n175), .Y(n149) );
  INVX1 U1380 ( .A(count[1]), .Y(n254) );
  INVX1 U1381 ( .A(n247), .Y(n246) );
  INVX1 U1382 ( .A(count[3]), .Y(n255) );
  OAI2BB1X1 U1383 ( .A0N(N327), .A1N(n974), .B0(n195), .Y(n748) );
  INVX1 U1384 ( .A(n936), .Y(n939) );
  INVX1 U1385 ( .A(n936), .Y(n938) );
  NOR2X1 U1386 ( .A(n1289), .B(n1288), .Y(n1290) );
  NAND4BXL U1387 ( .AN(n1287), .B(n856), .C(n1286), .D(n1285), .Y(n1289) );
  INVX1 U1388 ( .A(n259), .Y(n754) );
  AOI22X1 U1389 ( .A0(n969), .A1(count[8]), .B0(N278), .B1(n950), .Y(n259) );
  INVX1 U1390 ( .A(n260), .Y(n755) );
  AOI22X1 U1391 ( .A0(n969), .A1(count[7]), .B0(N277), .B1(n950), .Y(n260) );
  INVX1 U1392 ( .A(n261), .Y(n756) );
  AOI22X1 U1393 ( .A0(n969), .A1(count[6]), .B0(N276), .B1(n950), .Y(n261) );
  INVX1 U1394 ( .A(n262), .Y(n757) );
  AOI22X1 U1395 ( .A0(n969), .A1(count[5]), .B0(N275), .B1(n950), .Y(n262) );
  INVX1 U1396 ( .A(n263), .Y(n758) );
  AOI22X1 U1397 ( .A0(n969), .A1(count[4]), .B0(N274), .B1(n950), .Y(n263) );
  INVX1 U1398 ( .A(n264), .Y(n760) );
  AOI22X1 U1399 ( .A0(n969), .A1(count[2]), .B0(N272), .B1(n950), .Y(n264) );
  NAND2X1 U1400 ( .A(n106), .B(n1150), .Y(n1156) );
  OAI2BB2X1 U1401 ( .B0(n967), .B1(n255), .A0N(N273), .A1N(n950), .Y(n759) );
  OAI2BB2X1 U1402 ( .B0(n967), .B1(n254), .A0N(N271), .A1N(n950), .Y(n761) );
  NAND3X1 U1403 ( .A(count[1]), .B(n952), .C(n268), .Y(n1274) );
  INVX1 U1404 ( .A(n971), .Y(n973) );
  INVX1 U1405 ( .A(n971), .Y(n974) );
  OAI21XL U1406 ( .A0(n1149), .A1(n1148), .B0(N327), .Y(n72) );
  MXI2X1 U1407 ( .A(n142), .B(n1129), .S0(n1300), .Y(n1131) );
  NOR3X1 U1408 ( .A(n1128), .B(n1127), .C(n1126), .Y(n1129) );
  NAND2X1 U1409 ( .A(n1341), .B(n1332), .Y(n1127) );
  MX2X1 U1410 ( .A(n922), .B(n921), .S0(error_number[2]), .Y(N666) );
  MX4X1 U1411 ( .A(aadd1[7]), .B(aadd2[7]), .C(aadd3[7]), .D(aadd4[7]), .S0(
        n934), .S1(n938), .Y(n922) );
  MX4X1 U1412 ( .A(aadd5[7]), .B(aadd6[7]), .C(aadd7[7]), .D(aadd8[7]), .S0(
        n934), .S1(n938), .Y(n921) );
  MX2X1 U1413 ( .A(n930), .B(n929), .S0(error_number[2]), .Y(N662) );
  MX4X1 U1414 ( .A(aadd1[11]), .B(aadd2[11]), .C(aadd3[11]), .D(aadd4[11]), 
        .S0(n935), .S1(n939), .Y(n930) );
  MX4X1 U1415 ( .A(aadd5[11]), .B(aadd6[11]), .C(aadd7[11]), .D(aadd8[11]), 
        .S0(n935), .S1(n939), .Y(n929) );
  MX2X1 U1416 ( .A(n899), .B(n1311), .S0(n863), .Y(n1364) );
  AOI22X1 U1417 ( .A0(err_count[5]), .A1(n951), .B0(N668), .B1(n868), .Y(n80)
         );
  MX2X1 U1418 ( .A(n918), .B(n917), .S0(N258), .Y(N668) );
  MX4X1 U1419 ( .A(aadd1[5]), .B(aadd2[5]), .C(aadd3[5]), .D(aadd4[5]), .S0(
        n934), .S1(n938), .Y(n918) );
  MX2X1 U1420 ( .A(n932), .B(n931), .S0(error_number[2]), .Y(N661) );
  MX4X1 U1421 ( .A(aadd1[12]), .B(aadd2[12]), .C(aadd3[12]), .D(aadd4[12]), 
        .S0(n935), .S1(n939), .Y(n932) );
  AOI22X1 U1422 ( .A0(\add_587/carry[5] ), .A1(n951), .B0(N669), .B1(n868), 
        .Y(n93) );
  MX2X1 U1423 ( .A(n916), .B(n915), .S0(N258), .Y(N669) );
  MX4X1 U1424 ( .A(aadd1[4]), .B(aadd2[4]), .C(aadd3[4]), .D(aadd4[4]), .S0(
        n934), .S1(n938), .Y(n916) );
  AOI22X1 U1425 ( .A0(err_count[6]), .A1(n951), .B0(N667), .B1(n868), .Y(n94)
         );
  MX2X1 U1426 ( .A(n920), .B(n919), .S0(error_number[2]), .Y(N667) );
  MX4X1 U1427 ( .A(aadd1[6]), .B(aadd2[6]), .C(aadd3[6]), .D(aadd4[6]), .S0(
        n934), .S1(n938), .Y(n920) );
  NOR2X1 U1428 ( .A(n1281), .B(n1114), .Y(n1115) );
  NOR2X1 U1429 ( .A(n1288), .B(n1141), .Y(n1142) );
  NOR3X1 U1430 ( .A(sigma12[11]), .B(n1295), .C(n1296), .Y(n1134) );
  MX2X1 U1431 ( .A(n926), .B(n925), .S0(error_number[2]), .Y(N664) );
  MX4X1 U1432 ( .A(aadd1[9]), .B(aadd2[9]), .C(aadd3[9]), .D(aadd4[9]), .S0(
        n935), .S1(n939), .Y(n926) );
  MX4X1 U1433 ( .A(aadd5[9]), .B(aadd6[9]), .C(aadd7[9]), .D(aadd8[9]), .S0(
        n935), .S1(n939), .Y(n925) );
  MX2X1 U1434 ( .A(n928), .B(n927), .S0(error_number[2]), .Y(N663) );
  MX4X1 U1435 ( .A(aadd1[10]), .B(aadd2[10]), .C(aadd3[10]), .D(aadd4[10]), 
        .S0(n935), .S1(n939), .Y(n928) );
  MX4X1 U1436 ( .A(aadd5[10]), .B(aadd6[10]), .C(aadd7[10]), .D(aadd8[10]), 
        .S0(n935), .S1(n939), .Y(n927) );
  MX2X1 U1437 ( .A(n924), .B(n923), .S0(error_number[2]), .Y(N665) );
  MX4X1 U1438 ( .A(aadd1[8]), .B(aadd2[8]), .C(aadd3[8]), .D(aadd4[8]), .S0(
        n935), .S1(n939), .Y(n924) );
  MX4X1 U1439 ( .A(aadd5[8]), .B(aadd6[8]), .C(aadd7[8]), .D(aadd8[8]), .S0(
        n935), .S1(n939), .Y(n923) );
  NOR4X2 U1440 ( .A(n977), .B(e_sum_r[2]), .C(e_sum_r[3]), .D(e_sum_r[1]), .Y(
        n1107) );
  OAI22X1 U1441 ( .A0(n556), .A1(n116), .B0(n88), .B1(n117), .Y(n680) );
  OAI22X1 U1442 ( .A0(n558), .A1(n116), .B0(n90), .B1(n117), .Y(n682) );
  OAI22X1 U1443 ( .A0(n569), .A1(n121), .B0(n88), .B1(n122), .Y(n693) );
  OAI22X1 U1444 ( .A0(n571), .A1(n121), .B0(n90), .B1(n122), .Y(n695) );
  NAND3BX1 U1445 ( .AN(n235), .B(n597), .C(n820), .Y(n146) );
  NOR3X1 U1446 ( .A(sigma10[6]), .B(sigma10[4]), .C(sigma10[5]), .Y(n1002) );
  OAI2BB2X1 U1447 ( .B0(n1156), .B1(n84), .A0N(n949), .A1N(aadd1[1]), .Y(n644)
         );
  NAND3X1 U1448 ( .A(n974), .B(n951), .C(start_aadd), .Y(n152) );
  INVX1 U1449 ( .A(sigma8[6]), .Y(n1027) );
  NOR2X1 U1450 ( .A(sigma8[0]), .B(sigma8[1]), .Y(n1029) );
  NOR2X1 U1451 ( .A(sigma8[2]), .B(sigma8[3]), .Y(n1028) );
  OAI2BB2X1 U1452 ( .B0(n1156), .B1(n92), .A0N(n949), .A1N(aadd1[2]), .Y(n637)
         );
  OAI22X1 U1453 ( .A0(n485), .A1(n867), .B0(n80), .B1(n81), .Y(n609) );
  OAI22X1 U1454 ( .A0(n488), .A1(n79), .B0(n85), .B1(n81), .Y(n612) );
  OAI22X1 U1455 ( .A0(n496), .A1(n79), .B0(n93), .B1(n81), .Y(n620) );
  OAI22X1 U1456 ( .A0(n497), .A1(n867), .B0(n94), .B1(n81), .Y(n621) );
  OAI22X1 U1457 ( .A0(n498), .A1(n98), .B0(n80), .B1(n99), .Y(n622) );
  OAI22X1 U1458 ( .A0(n501), .A1(n98), .B0(n85), .B1(n99), .Y(n625) );
  OAI22X1 U1459 ( .A0(n509), .A1(n98), .B0(n93), .B1(n99), .Y(n633) );
  OAI22X1 U1460 ( .A0(n510), .A1(n860), .B0(n94), .B1(n99), .Y(n634) );
  OAI22X1 U1461 ( .A0(n511), .A1(n1504), .B0(n94), .B1(n1629), .Y(n635) );
  OAI22X1 U1462 ( .A0(n512), .A1(n1504), .B0(n93), .B1(n1629), .Y(n636) );
  OAI22X1 U1463 ( .A0(n519), .A1(n1504), .B0(n85), .B1(n1629), .Y(n643) );
  OAI22X1 U1464 ( .A0(n522), .A1(n1504), .B0(n80), .B1(n1629), .Y(n646) );
  OAI22X1 U1465 ( .A0(n524), .A1(n107), .B0(n94), .B1(n108), .Y(n648) );
  OAI22X1 U1466 ( .A0(n525), .A1(n866), .B0(n93), .B1(n108), .Y(n649) );
  OAI22X1 U1467 ( .A0(n532), .A1(n107), .B0(n85), .B1(n108), .Y(n656) );
  OAI22X1 U1468 ( .A0(n535), .A1(n107), .B0(n80), .B1(n108), .Y(n659) );
  OAI22X1 U1469 ( .A0(n537), .A1(n111), .B0(n94), .B1(n112), .Y(n661) );
  OAI22X1 U1470 ( .A0(n538), .A1(n111), .B0(n93), .B1(n112), .Y(n662) );
  OAI22X1 U1471 ( .A0(n545), .A1(n111), .B0(n85), .B1(n112), .Y(n669) );
  OAI22X1 U1472 ( .A0(n548), .A1(n111), .B0(n80), .B1(n112), .Y(n672) );
  OAI22X1 U1473 ( .A0(n550), .A1(n865), .B0(n80), .B1(n117), .Y(n674) );
  OAI22X1 U1474 ( .A0(n553), .A1(n116), .B0(n85), .B1(n117), .Y(n677) );
  OAI22X1 U1475 ( .A0(n561), .A1(n116), .B0(n93), .B1(n117), .Y(n685) );
  OAI22X1 U1476 ( .A0(n562), .A1(n865), .B0(n94), .B1(n117), .Y(n686) );
  OAI22X1 U1477 ( .A0(n563), .A1(n121), .B0(n80), .B1(n122), .Y(n687) );
  OAI22X1 U1478 ( .A0(n566), .A1(n121), .B0(n85), .B1(n122), .Y(n690) );
  OAI22X1 U1479 ( .A0(n574), .A1(n121), .B0(n93), .B1(n122), .Y(n698) );
  OAI22X1 U1480 ( .A0(n575), .A1(n121), .B0(n94), .B1(n122), .Y(n699) );
  OAI22X1 U1481 ( .A0(n576), .A1(n864), .B0(n80), .B1(n125), .Y(n700) );
  OAI22X1 U1482 ( .A0(n579), .A1(n124), .B0(n85), .B1(n125), .Y(n703) );
  OAI22X1 U1483 ( .A0(n587), .A1(n124), .B0(n93), .B1(n125), .Y(n711) );
  OAI22X1 U1484 ( .A0(n588), .A1(n864), .B0(n94), .B1(n125), .Y(n712) );
  NOR2X1 U1485 ( .A(sigma2[0]), .B(sigma2[1]), .Y(n1013) );
  NOR2X1 U1486 ( .A(sigma2[2]), .B(sigma2[3]), .Y(n1012) );
  NOR2X1 U1487 ( .A(sigma16[6]), .B(sigma16[8]), .Y(n1091) );
  NOR2X1 U1488 ( .A(sigma16[9]), .B(sigma16[12]), .Y(n1089) );
  NOR2X1 U1489 ( .A(sigma13[6]), .B(sigma13[8]), .Y(n1085) );
  NOR2X1 U1490 ( .A(sigma13[9]), .B(sigma13[12]), .Y(n1083) );
  NOR2X1 U1491 ( .A(sigma3[0]), .B(sigma3[1]), .Y(n1007) );
  INVX1 U1492 ( .A(sigma3[6]), .Y(n1005) );
  NOR2X1 U1493 ( .A(sigma3[2]), .B(sigma3[3]), .Y(n1006) );
  NOR2X1 U1494 ( .A(n605), .B(n765), .Y(n199) );
  NOR2X1 U1495 ( .A(sigma12[6]), .B(sigma12[8]), .Y(n1019) );
  INVX1 U1496 ( .A(sigma12[7]), .Y(n1018) );
  NOR2X1 U1497 ( .A(sigma12[9]), .B(sigma12[12]), .Y(n1017) );
  NOR3X1 U1498 ( .A(sigma5[6]), .B(sigma5[4]), .C(sigma5[5]), .Y(n1079) );
  NOR3X1 U1499 ( .A(sigma5[9]), .B(sigma5[7]), .C(sigma5[8]), .Y(n1078) );
  NOR3X1 U1500 ( .A(sigma5[12]), .B(sigma5[10]), .C(sigma5[11]), .Y(n1077) );
  XOR3X2 U1501 ( .A(n940), .B(n1458), .C(n1420), .Y(n901) );
  INVX1 U1502 ( .A(e_sum_r[0]), .Y(n1359) );
  OAI2BB2X1 U1503 ( .B0(n1156), .B1(n91), .A0N(n949), .A1N(aadd1[0]), .Y(n638)
         );
  OAI2BB2X1 U1504 ( .B0(n1156), .B1(n83), .A0N(n949), .A1N(aadd1[3]), .Y(n645)
         );
  OAI22X1 U1505 ( .A0(n196), .A1(n976), .B0(N256), .B1(n152), .Y(n737) );
  NOR3X1 U1506 ( .A(sigma6[9]), .B(sigma6[7]), .C(sigma6[8]), .Y(n1070) );
  OAI2BB1X1 U1507 ( .A0N(n140), .A1N(n141), .B0(n974), .Y(n91) );
  AOI21X1 U1508 ( .A0(n765), .A1(n142), .B0(n143), .Y(n140) );
  MX2X1 U1509 ( .A(n908), .B(n907), .S0(error_number[2]), .Y(N673) );
  NOR3X1 U1510 ( .A(sigma8[12]), .B(sigma8[10]), .C(sigma8[11]), .Y(n1030) );
  NOR3X1 U1511 ( .A(sigma8[9]), .B(sigma8[7]), .C(sigma8[8]), .Y(n1031) );
  NOR2X1 U1512 ( .A(n1656), .B(sigma14[0]), .Y(n1135) );
  NOR2X1 U1513 ( .A(n1649), .B(sigma11[8]), .Y(n1065) );
  NOR2X1 U1514 ( .A(sigma7[4]), .B(sigma7[5]), .Y(n993) );
  NOR2X1 U1515 ( .A(sigma4[4]), .B(sigma4[5]), .Y(n987) );
  OAI22X1 U1516 ( .A0(n118), .A1(n83), .B0(n551), .B1(n865), .Y(n675) );
  OAI22X1 U1517 ( .A0(n118), .A1(n91), .B0(n559), .B1(n865), .Y(n683) );
  OAI22X1 U1518 ( .A0(n123), .A1(n83), .B0(n564), .B1(n858), .Y(n688) );
  OAI22X1 U1519 ( .A0(n123), .A1(n91), .B0(n572), .B1(n858), .Y(n696) );
  OAI22X1 U1520 ( .A0(n82), .A1(n83), .B0(n486), .B1(n867), .Y(n610) );
  OAI22X1 U1521 ( .A0(n82), .A1(n91), .B0(n494), .B1(n867), .Y(n618) );
  OAI22X1 U1522 ( .A0(n100), .A1(n83), .B0(n499), .B1(n860), .Y(n623) );
  OAI22X1 U1523 ( .A0(n100), .A1(n91), .B0(n507), .B1(n860), .Y(n631) );
  OAI22X1 U1524 ( .A0(n109), .A1(n91), .B0(n527), .B1(n866), .Y(n651) );
  OAI22X1 U1525 ( .A0(n109), .A1(n83), .B0(n534), .B1(n866), .Y(n658) );
  OAI22X1 U1526 ( .A0(n113), .A1(n91), .B0(n540), .B1(n859), .Y(n664) );
  OAI22X1 U1527 ( .A0(n113), .A1(n83), .B0(n547), .B1(n859), .Y(n671) );
  OAI22X1 U1528 ( .A0(n129), .A1(n83), .B0(n577), .B1(n864), .Y(n701) );
  OAI22X1 U1529 ( .A0(n129), .A1(n91), .B0(n585), .B1(n864), .Y(n709) );
  NAND3X1 U1530 ( .A(n210), .B(n899), .C(n764), .Y(n200) );
  NAND4X2 U1531 ( .A(n984), .B(n985), .C(n983), .D(n982), .Y(n1106) );
  NOR2X1 U1532 ( .A(n979), .B(n589), .Y(n985) );
  NAND4X1 U1533 ( .A(n1062), .B(n1061), .C(n1060), .D(n1059), .Y(n1130) );
  NOR3XL U1534 ( .A(sigma9[4]), .B(n1648), .C(n1647), .Y(n1060) );
  NOR3XL U1535 ( .A(sigma9[1]), .B(sigma9[0]), .C(sigma9[2]), .Y(n1059) );
  NOR3X1 U1536 ( .A(sigma2[8]), .B(sigma2[9]), .C(sigma2[7]), .Y(n1033) );
  OAI21XL U1537 ( .A0(n1300), .A1(n149), .B0(n968), .Y(n1162) );
  NAND4X1 U1538 ( .A(n1042), .B(n1041), .C(n1040), .D(n1039), .Y(n1049) );
  NOR2XL U1539 ( .A(sigma13[0]), .B(sigma14[12]), .Y(n1042) );
  AND2X2 U1540 ( .A(n214), .B(n603), .Y(n138) );
  NAND3BX1 U1541 ( .AN(n206), .B(n593), .C(n821), .Y(n77) );
  INVX1 U1542 ( .A(sigma16[10]), .Y(n1050) );
  NOR2X1 U1543 ( .A(sigma15[1]), .B(sigma15[0]), .Y(n1052) );
  NAND2X1 U1544 ( .A(n604), .B(n210), .Y(n165) );
  OAI21XL U1545 ( .A0(n1300), .A1(n138), .B0(n968), .Y(n1159) );
  OAI2BB2X1 U1546 ( .B0(n589), .B1(n902), .A0N(N817), .A1N(n1505), .Y(n723) );
  NAND2X1 U1547 ( .A(n1112), .B(n1111), .Y(n1280) );
  NAND2X1 U1548 ( .A(n1138), .B(n1137), .Y(n1287) );
  NOR2X1 U1549 ( .A(sigma15[3]), .B(sigma15[2]), .Y(n1053) );
  XNOR3X2 U1550 ( .A(n1400), .B(n1399), .C(n1398), .Y(n1401) );
  NOR2X1 U1551 ( .A(sigma14[9]), .B(sigma14[8]), .Y(n1023) );
  NOR2X1 U1552 ( .A(sigma15[9]), .B(sigma15[8]), .Y(n1021) );
  NOR2X1 U1553 ( .A(sigma14[7]), .B(sigma14[6]), .Y(n1022) );
  NOR2X1 U1554 ( .A(sigma15[7]), .B(sigma15[6]), .Y(n1020) );
  NOR2X1 U1555 ( .A(sigma7[0]), .B(sigma7[1]), .Y(n995) );
  NOR2X1 U1556 ( .A(sigma4[0]), .B(sigma4[1]), .Y(n989) );
  OAI2BB2X1 U1557 ( .B0(n590), .B1(n902), .A0N(N811), .A1N(n1505), .Y(n729) );
  OAI2BB2X1 U1558 ( .B0(n591), .B1(n902), .A0N(N810), .A1N(n1505), .Y(n730) );
  OAI2BB2X1 U1559 ( .B0(n592), .B1(n902), .A0N(n592), .A1N(n1505), .Y(n731) );
  NOR2X1 U1560 ( .A(sigma7[2]), .B(sigma7[3]), .Y(n994) );
  NOR2X1 U1561 ( .A(sigma4[2]), .B(sigma4[3]), .Y(n988) );
  OR2X2 U1562 ( .A(sigma11[10]), .B(sigma11[0]), .Y(n1302) );
  NOR2X1 U1563 ( .A(sigma12[1]), .B(sigma12[3]), .Y(n1016) );
  NOR2X1 U1564 ( .A(n1654), .B(sigma12[5]), .Y(n1014) );
  NOR2X1 U1565 ( .A(sigma16[1]), .B(sigma16[3]), .Y(n1094) );
  NOR2X1 U1566 ( .A(sigma16[4]), .B(sigma16[5]), .Y(n1092) );
  NOR2X1 U1567 ( .A(sigma13[1]), .B(sigma13[3]), .Y(n1088) );
  INVX1 U1568 ( .A(sigma13[2]), .Y(n1087) );
  NOR2X1 U1569 ( .A(n1653), .B(n1651), .Y(n1068) );
  NOR2X1 U1570 ( .A(n1650), .B(sigma11[5]), .Y(n1066) );
  NAND2X1 U1571 ( .A(n603), .B(n1397), .Y(n1383) );
  AND4X2 U1572 ( .A(n165), .B(n200), .C(n201), .D(n202), .Y(n130) );
  NOR2X1 U1573 ( .A(n602), .B(n138), .Y(n201) );
  AND4X2 U1574 ( .A(n135), .B(n147), .C(n175), .D(n813), .Y(n202) );
  MX4X1 U1575 ( .A(aadd1[1]), .B(aadd2[1]), .C(aadd3[1]), .D(aadd4[1]), .S0(
        error_number[0]), .S1(error_number[1]), .Y(n910) );
  MX4X1 U1576 ( .A(aadd1[2]), .B(aadd2[2]), .C(aadd3[2]), .D(aadd4[2]), .S0(
        error_number[0]), .S1(error_number[1]), .Y(n912) );
  AOI2BB2X1 U1577 ( .B0(n600), .B1(n1161), .A0N(n857), .A1N(n1332), .Y(n719)
         );
  OAI21XL U1578 ( .A0(n1300), .A1(n172), .B0(n968), .Y(n1161) );
  AOI2BB2X1 U1579 ( .B0(n602), .B1(n1163), .A0N(n857), .A1N(n1343), .Y(n721)
         );
  OAI21XL U1580 ( .A0(n1300), .A1(n813), .B0(n968), .Y(n1163) );
  NAND2X1 U1581 ( .A(n1044), .B(n1043), .Y(n1048) );
  NOR2XL U1582 ( .A(sigma12[10]), .B(sigma12[0]), .Y(n1044) );
  NOR2XL U1583 ( .A(sigma13[11]), .B(sigma13[10]), .Y(n1043) );
  MX4X1 U1584 ( .A(aadd5[1]), .B(aadd6[1]), .C(aadd7[1]), .D(aadd8[1]), .S0(
        error_number[0]), .S1(error_number[1]), .Y(n909) );
  MX4X1 U1585 ( .A(aadd5[2]), .B(aadd6[2]), .C(aadd7[2]), .D(aadd8[2]), .S0(
        error_number[0]), .S1(error_number[1]), .Y(n911) );
  OAI21XL U1586 ( .A0(n1300), .A1(n160), .B0(n968), .Y(n1157) );
  OAI21XL U1587 ( .A0(n1300), .A1(n212), .B0(n968), .Y(n1283) );
  NAND4BXL U1588 ( .AN(n1280), .B(n856), .C(n1279), .D(n1278), .Y(n1282) );
  AOI21X1 U1589 ( .A0(n596), .A1(n1294), .B0(n1293), .Y(n740) );
  OAI21XL U1590 ( .A0(n1300), .A1(n211), .B0(n968), .Y(n1294) );
  AOI21X1 U1591 ( .A0(n598), .A1(n1304), .B0(n1303), .Y(n742) );
  OAI21XL U1592 ( .A0(n1300), .A1(n145), .B0(n968), .Y(n1304) );
  INVX1 U1593 ( .A(error_number[3]), .Y(n1277) );
  INVX1 U1594 ( .A(sigma15[12]), .Y(n1279) );
  AOI21X1 U1595 ( .A0(n971), .A1(e_sum_r[3]), .B0(n1475), .Y(n1476) );
  INVX1 U1596 ( .A(n1488), .Y(n1475) );
  INVX1 U1597 ( .A(n181), .Y(n724) );
  INVX1 U1598 ( .A(n183), .Y(n725) );
  INVX1 U1599 ( .A(n184), .Y(n726) );
  INVX1 U1600 ( .A(n185), .Y(n727) );
  INVX1 U1601 ( .A(n186), .Y(n728) );
  NOR3X1 U1602 ( .A(sigma4[9]), .B(sigma4[7]), .C(sigma4[8]), .Y(n991) );
  NOR3X1 U1603 ( .A(sigma4[12]), .B(sigma4[10]), .C(sigma4[11]), .Y(n990) );
  MX2X1 U1604 ( .A(n914), .B(n913), .S0(N258), .Y(N670) );
  MX4X1 U1605 ( .A(aadd1[3]), .B(aadd2[3]), .C(aadd3[3]), .D(aadd4[3]), .S0(
        n934), .S1(n938), .Y(n914) );
  INVX1 U1606 ( .A(sigma2[5]), .Y(n1010) );
  INVX1 U1607 ( .A(sigma7[6]), .Y(n992) );
  INVX1 U1608 ( .A(sigma4[6]), .Y(n986) );
  OAI32X1 U1609 ( .A0(n152), .A1(N258), .A2(n153), .B0(n154), .B1(n115), .Y(
        n713) );
  NOR2X1 U1610 ( .A(n153), .B(n155), .Y(n154) );
  INVX1 U1611 ( .A(n902), .Y(n182) );
  INVX1 U1612 ( .A(N1190), .Y(n975) );
  INVX1 U1613 ( .A(n156), .Y(n714) );
  INVX1 U1614 ( .A(n152), .Y(n157) );
  NOR3BX1 U1615 ( .AN(count[6]), .B(count[0]), .C(count[2]), .Y(n268) );
  NOR3X1 U1616 ( .A(count[7]), .B(count[9]), .C(count[8]), .Y(n256) );
  INVX1 U1617 ( .A(n265), .Y(n762) );
  AOI22X1 U1618 ( .A0(n971), .A1(count[0]), .B0(N270), .B1(n950), .Y(n265) );
  OAI2BB1X1 U1619 ( .A0N(Uin[0]), .A1N(n247), .B0(n249), .Y(n752) );
  NAND4BXL U1620 ( .AN(count[0]), .B(n250), .C(n246), .D(n251), .Y(n249) );
  MXI2X1 U1621 ( .A(n1265), .B(n1266), .S0(n953), .Y(n1520) );
  INVX1 U1622 ( .A(err_loc8[12]), .Y(n1265) );
  MXI2X1 U1623 ( .A(n1203), .B(n1204), .S0(n959), .Y(n1583) );
  INVX1 U1624 ( .A(err_loc8[5]), .Y(n1203) );
  MXI2X1 U1625 ( .A(n1276), .B(n1275), .S0(n954), .Y(N449) );
  INVX1 U1626 ( .A(sel_ch), .Y(n1276) );
  MXI2X1 U1627 ( .A(n1194), .B(n1195), .S0(n960), .Y(n1592) );
  INVX1 U1628 ( .A(err_loc8[4]), .Y(n1194) );
  MXI2X1 U1629 ( .A(n1176), .B(n1177), .S0(n961), .Y(n1610) );
  INVX1 U1630 ( .A(err_loc8[2]), .Y(n1176) );
  MXI2X1 U1631 ( .A(n1185), .B(n1186), .S0(n961), .Y(n1601) );
  INVX1 U1632 ( .A(err_loc8[3]), .Y(n1185) );
  MXI2X1 U1633 ( .A(n1238), .B(n1239), .S0(n956), .Y(n1547) );
  INVX1 U1634 ( .A(err_loc8[9]), .Y(n1238) );
  MXI2X1 U1635 ( .A(n1229), .B(n1230), .S0(n956), .Y(n1556) );
  INVX1 U1636 ( .A(err_loc8[8]), .Y(n1229) );
  MXI2X1 U1637 ( .A(n1212), .B(n1213), .S0(n958), .Y(n1574) );
  INVX1 U1638 ( .A(err_loc8[6]), .Y(n1212) );
  MXI2X1 U1639 ( .A(n1247), .B(n1248), .S0(n955), .Y(n1538) );
  INVX1 U1640 ( .A(err_loc8[10]), .Y(n1247) );
  MXI2X1 U1641 ( .A(n1256), .B(n1257), .S0(n954), .Y(n1529) );
  INVX1 U1642 ( .A(err_loc8[11]), .Y(n1256) );
  MXI2X1 U1643 ( .A(n1175), .B(n1174), .S0(n961), .Y(n1612) );
  INVX1 U1644 ( .A(err_loc0[1]), .Y(n1174) );
  MXI2X1 U1645 ( .A(n1184), .B(n1183), .S0(n960), .Y(n1603) );
  INVX1 U1646 ( .A(err_loc0[2]), .Y(n1183) );
  MXI2X1 U1647 ( .A(n1193), .B(n1192), .S0(n960), .Y(n1594) );
  INVX1 U1648 ( .A(err_loc0[3]), .Y(n1192) );
  MXI2X1 U1649 ( .A(n1202), .B(n1201), .S0(n959), .Y(n1585) );
  INVX1 U1650 ( .A(err_loc0[4]), .Y(n1201) );
  MXI2X1 U1651 ( .A(n1211), .B(n1210), .S0(n958), .Y(n1576) );
  INVX1 U1652 ( .A(err_loc0[5]), .Y(n1210) );
  MXI2X1 U1653 ( .A(n1220), .B(n1219), .S0(n957), .Y(n1567) );
  INVX1 U1654 ( .A(err_loc0[6]), .Y(n1219) );
  MXI2X1 U1655 ( .A(n1228), .B(n1227), .S0(n957), .Y(n1558) );
  INVX1 U1656 ( .A(err_loc0[7]), .Y(n1227) );
  MXI2X1 U1657 ( .A(n1237), .B(n1236), .S0(n956), .Y(n1549) );
  INVX1 U1658 ( .A(err_loc0[8]), .Y(n1236) );
  MXI2X1 U1659 ( .A(n1246), .B(n1245), .S0(n955), .Y(n1540) );
  INVX1 U1660 ( .A(err_loc0[9]), .Y(n1245) );
  MXI2X1 U1661 ( .A(n1255), .B(n1254), .S0(n954), .Y(n1531) );
  INVX1 U1662 ( .A(err_loc0[10]), .Y(n1254) );
  MXI2X1 U1663 ( .A(n1264), .B(n1263), .S0(n953), .Y(n1522) );
  INVX1 U1664 ( .A(err_loc0[11]), .Y(n1263) );
  MXI2X1 U1665 ( .A(n1273), .B(n1272), .S0(n953), .Y(n1513) );
  INVX1 U1666 ( .A(err_loc0[12]), .Y(n1272) );
  AOI22X1 U1667 ( .A0(n597), .A1(n1299), .B0(n1298), .B1(n1297), .Y(n741) );
  NOR2X1 U1668 ( .A(n1295), .B(n857), .Y(n1298) );
  NAND2X1 U1669 ( .A(n1307), .B(n1306), .Y(n743) );
  INVX1 U1670 ( .A(start_aadd), .Y(n195) );
  OAI2BB1X1 U1671 ( .A0N(n135), .A1N(n1309), .B0(n973), .Y(n1160) );
  AOI22X1 U1672 ( .A0(n593), .A1(n1155), .B0(n1154), .B1(n1153), .Y(n608) );
  NOR2X1 U1673 ( .A(n1151), .B(n857), .Y(n1154) );
  MX4X1 U1674 ( .A(aadd1[0]), .B(aadd2[0]), .C(aadd3[0]), .D(aadd4[0]), .S0(
        error_number[0]), .S1(error_number[1]), .Y(n908) );
  AOI2BB2X1 U1675 ( .B0(n604), .B1(n1158), .A0N(n857), .A1N(n1311), .Y(n716)
         );
  OAI2BB1X1 U1676 ( .A0N(n165), .A1N(n875), .B0(n973), .Y(n1158) );
  MX4X1 U1677 ( .A(aadd5[3]), .B(aadd6[3]), .C(aadd7[3]), .D(aadd8[3]), .S0(
        n934), .S1(n938), .Y(n913) );
  MX4X1 U1678 ( .A(aadd5[0]), .B(aadd6[0]), .C(aadd7[0]), .D(aadd8[0]), .S0(
        error_number[0]), .S1(error_number[1]), .Y(n907) );
  MX4X1 U1679 ( .A(aadd5[5]), .B(aadd6[5]), .C(aadd7[5]), .D(aadd8[5]), .S0(
        n934), .S1(n938), .Y(n917) );
  MX4X1 U1680 ( .A(aadd5[12]), .B(aadd6[12]), .C(aadd7[12]), .D(aadd8[12]), 
        .S0(n935), .S1(n939), .Y(n931) );
  MX4X1 U1681 ( .A(aadd5[4]), .B(aadd6[4]), .C(aadd7[4]), .D(aadd8[4]), .S0(
        n934), .S1(n938), .Y(n915) );
  MX4X1 U1682 ( .A(aadd5[6]), .B(aadd6[6]), .C(aadd7[6]), .D(aadd8[6]), .S0(
        n934), .S1(n938), .Y(n919) );
  NAND4X1 U1683 ( .A(count[9]), .B(count[8]), .C(count[7]), .D(count[5]), .Y(
        n267) );
  NAND4BXL U1684 ( .AN(n952), .B(n268), .C(count[3]), .D(n254), .Y(n266) );
  OAI31X1 U1685 ( .A0(n252), .A1(N266), .A2(n250), .B0(n973), .Y(n247) );
  NAND2X1 U1686 ( .A(n251), .B(n248), .Y(n252) );
  BUFX3 U1687 ( .A(count[4]), .Y(n952) );
  NOR2X1 U1688 ( .A(n606), .B(n246), .Y(n749) );
  MX2X1 U1689 ( .A(err_loc0[0]), .B(Lout[0]), .S0(n964), .Y(n1620) );
  MX2X1 U1690 ( .A(err_loc0[1]), .B(Lout[1]), .S0(n964), .Y(n1611) );
  MX2X1 U1691 ( .A(err_loc0[2]), .B(Lout[2]), .S0(n964), .Y(n1602) );
  MX2X1 U1692 ( .A(err_loc0[3]), .B(Lout[3]), .S0(n963), .Y(n1593) );
  MX2X1 U1693 ( .A(err_loc0[4]), .B(Lout[4]), .S0(n963), .Y(n1584) );
  MX2X1 U1694 ( .A(err_loc0[5]), .B(Lout[5]), .S0(n963), .Y(n1575) );
  MX2X1 U1695 ( .A(err_loc0[6]), .B(Lout[6]), .S0(n964), .Y(n1566) );
  MX2X1 U1696 ( .A(err_loc0[7]), .B(Lout[7]), .S0(n964), .Y(n1557) );
  MX2X1 U1697 ( .A(err_loc0[8]), .B(Lout[8]), .S0(n963), .Y(n1548) );
  MX2X1 U1698 ( .A(err_loc0[9]), .B(Lout[9]), .S0(n964), .Y(n1539) );
  MX2X1 U1699 ( .A(err_loc0[10]), .B(Lout[10]), .S0(n964), .Y(n1530) );
  MX2X1 U1700 ( .A(err_loc0[11]), .B(Lout[11]), .S0(n964), .Y(n1521) );
  MX2X1 U1701 ( .A(err_loc0[12]), .B(Lout[12]), .S0(n964), .Y(n1512) );
  OR2X2 U1702 ( .A(start_eu), .B(n246), .Y(n751) );
  OAI32X1 U1703 ( .A0(n247), .A1(count[0]), .A2(n248), .B0(n246), .B1(n607), 
        .Y(n750) );
  INVX1 U1704 ( .A(n257), .Y(n753) );
  AOI22X1 U1705 ( .A0(n971), .A1(count[9]), .B0(N279), .B1(n950), .Y(n257) );
  INVX1 U1706 ( .A(err_loc3[12]), .Y(n1270) );
  INVX1 U1707 ( .A(err_loc6[4]), .Y(n1196) );
  INVX1 U1708 ( .A(err_loc7[12]), .Y(n1266) );
  INVX1 U1709 ( .A(err_loc2[1]), .Y(n1173) );
  INVX1 U1710 ( .A(err_loc5[4]), .Y(n1197) );
  INVX1 U1711 ( .A(err_loc7[5]), .Y(n1204) );
  INVX1 U1712 ( .A(err_loc1[11]), .Y(n1264) );
  INVX1 U1713 ( .A(err_loc6[12]), .Y(n1267) );
  INVX1 U1714 ( .A(err_loc2[8]), .Y(n1235) );
  INVX1 U1715 ( .A(err_loc5[5]), .Y(n1206) );
  INVX1 U1716 ( .A(err_loc4[2]), .Y(n1180) );
  INVX1 U1717 ( .A(err_loc5[6]), .Y(n1215) );
  INVX1 U1718 ( .A(err_loc2[6]), .Y(n1218) );
  INVX1 U1719 ( .A(err_loc4[9]), .Y(n1242) );
  INVX1 U1720 ( .A(err_loc2[9]), .Y(n1244) );
  INVX1 U1721 ( .A(err_loc4[0]), .Y(n1166) );
  INVX1 U1722 ( .A(err_loc4[1]), .Y(n1171) );
  INVX1 U1723 ( .A(err_loc5[2]), .Y(n1179) );
  INVX1 U1724 ( .A(err_loc2[2]), .Y(n1182) );
  INVX1 U1725 ( .A(err_loc1[2]), .Y(n1184) );
  INVX1 U1726 ( .A(err_loc4[4]), .Y(n1198) );
  INVX1 U1727 ( .A(err_loc1[4]), .Y(n1202) );
  INVX1 U1728 ( .A(err_loc4[5]), .Y(n1207) );
  INVX1 U1729 ( .A(err_loc7[7]), .Y(n1221) );
  INVX1 U1730 ( .A(err_loc2[7]), .Y(n1226) );
  INVX1 U1731 ( .A(err_loc1[7]), .Y(n1228) );
  INVX1 U1732 ( .A(err_loc4[8]), .Y(n1233) );
  INVX1 U1733 ( .A(err_loc1[8]), .Y(n1237) );
  INVX1 U1734 ( .A(err_loc6[11]), .Y(n1258) );
  INVX1 U1735 ( .A(err_loc2[11]), .Y(n1262) );
  INVX1 U1736 ( .A(err_loc5[1]), .Y(n1170) );
  INVX1 U1737 ( .A(err_loc6[3]), .Y(n1187) );
  INVX1 U1738 ( .A(err_loc7[4]), .Y(n1195) );
  INVX1 U1739 ( .A(err_loc7[2]), .Y(n1177) );
  INVX1 U1740 ( .A(err_loc5[3]), .Y(n1188) );
  INVX1 U1741 ( .A(err_loc4[3]), .Y(n1189) );
  INVX1 U1742 ( .A(err_loc6[8]), .Y(n1231) );
  INVX1 U1743 ( .A(err_loc4[10]), .Y(n1251) );
  INVX1 U1744 ( .A(err_loc2[10]), .Y(n1253) );
  INVX1 U1745 ( .A(err_loc7[3]), .Y(n1186) );
  INVX1 U1746 ( .A(err_loc5[7]), .Y(n1223) );
  INVX1 U1747 ( .A(err_loc5[9]), .Y(n1241) );
  INVX1 U1748 ( .A(err_loc4[12]), .Y(n1269) );
  INVX1 U1749 ( .A(err_loc2[0]), .Y(n1168) );
  INVX1 U1750 ( .A(err_loc2[5]), .Y(n1209) );
  INVX1 U1751 ( .A(err_loc7[9]), .Y(n1239) );
  INVX1 U1752 ( .A(err_loc1[9]), .Y(n1246) );
  INVX1 U1753 ( .A(err_loc6[6]), .Y(n1214) );
  INVX1 U1754 ( .A(err_loc1[6]), .Y(n1220) );
  INVX1 U1755 ( .A(err_loc7[8]), .Y(n1230) );
  INVX1 U1756 ( .A(err_loc1[10]), .Y(n1255) );
  INVX1 U1757 ( .A(err_loc4[11]), .Y(n1260) );
  INVX1 U1758 ( .A(err_loc5[0]), .Y(n1165) );
  INVX1 U1759 ( .A(err_loc3[3]), .Y(n1190) );
  INVX1 U1760 ( .A(err_loc5[11]), .Y(n1259) );
  INVX1 U1761 ( .A(err_loc3[0]), .Y(n1167) );
  INVX1 U1762 ( .A(err_loc6[1]), .Y(n1169) );
  INVX1 U1763 ( .A(err_loc3[1]), .Y(n1172) );
  INVX1 U1764 ( .A(err_loc1[3]), .Y(n1193) );
  INVX1 U1765 ( .A(err_loc3[4]), .Y(n1199) );
  INVX1 U1766 ( .A(err_loc3[5]), .Y(n1208) );
  INVX1 U1767 ( .A(err_loc4[6]), .Y(n1216) );
  INVX1 U1768 ( .A(err_loc3[6]), .Y(n1217) );
  INVX1 U1769 ( .A(err_loc6[7]), .Y(n1222) );
  INVX1 U1770 ( .A(err_loc5[8]), .Y(n1232) );
  INVX1 U1771 ( .A(err_loc3[11]), .Y(n1261) );
  INVX1 U1772 ( .A(err_loc4[7]), .Y(n1224) );
  INVX1 U1773 ( .A(err_loc3[8]), .Y(n1234) );
  INVX1 U1774 ( .A(err_loc3[7]), .Y(n1225) );
  INVX1 U1775 ( .A(err_loc6[9]), .Y(n1240) );
  INVX1 U1776 ( .A(err_loc6[0]), .Y(n1164) );
  INVX1 U1777 ( .A(err_loc1[1]), .Y(n1175) );
  INVX1 U1778 ( .A(err_loc6[2]), .Y(n1178) );
  INVX1 U1779 ( .A(err_loc2[3]), .Y(n1191) );
  INVX1 U1780 ( .A(err_loc2[4]), .Y(n1200) );
  INVX1 U1781 ( .A(err_loc1[5]), .Y(n1211) );
  INVX1 U1782 ( .A(err_loc7[6]), .Y(n1213) );
  INVX1 U1783 ( .A(err_loc5[10]), .Y(n1250) );
  INVX1 U1784 ( .A(err_loc3[10]), .Y(n1252) );
  INVX1 U1785 ( .A(err_loc2[12]), .Y(n1271) );
  INVX1 U1786 ( .A(err_loc1[12]), .Y(n1273) );
  INVX1 U1787 ( .A(err_loc3[2]), .Y(n1181) );
  INVX1 U1788 ( .A(err_loc6[5]), .Y(n1205) );
  INVX1 U1789 ( .A(err_loc7[10]), .Y(n1248) );
  INVX1 U1790 ( .A(err_loc6[10]), .Y(n1249) );
  INVX1 U1791 ( .A(err_loc7[11]), .Y(n1257) );
  INVX1 U1792 ( .A(err_loc5[12]), .Y(n1268) );
  INVX1 U1793 ( .A(err_loc3[9]), .Y(n1243) );
  NOR4X1 U1794 ( .A(n286), .B(n287), .C(n288), .D(n289), .Y(error_finish) );
  NAND4X1 U1795 ( .A(n596), .B(n595), .C(n594), .D(n593), .Y(n286) );
  NAND4X1 U1796 ( .A(n599), .B(n605), .C(n598), .D(n597), .Y(n287) );
  NOR3X1 U1797 ( .A(n72), .B(n269), .C(n195), .Y(error_occur) );
  MXI2XL U1802 ( .A(n764), .B(n1310), .S0(n974), .Y(N1141) );
  NAND4BXL U1803 ( .AN(n765), .B(n874), .C(n142), .D(n973), .Y(n1306) );
  MXI2X1 U1804 ( .A(n1359), .B(n1358), .S0(n973), .Y(n1511) );
  NAND4X1 U1805 ( .A(n101), .B(n97), .C(n974), .D(n951), .Y(n194) );
  OAI22X1 U1806 ( .A0(n584), .A1(n124), .B0(n90), .B1(n125), .Y(n708) );
  OAI22X1 U1807 ( .A0(n493), .A1(n79), .B0(n90), .B1(n81), .Y(n617) );
  OAI22X1 U1808 ( .A0(n506), .A1(n98), .B0(n90), .B1(n99), .Y(n630) );
  OAI22X1 U1809 ( .A0(n515), .A1(n1504), .B0(n90), .B1(n949), .Y(n639) );
  OAI22X1 U1810 ( .A0(n528), .A1(n107), .B0(n90), .B1(n108), .Y(n652) );
  OAI22X1 U1811 ( .A0(n541), .A1(n111), .B0(n90), .B1(n112), .Y(n665) );
  OAI22X1 U1812 ( .A0(n492), .A1(n79), .B0(n89), .B1(n81), .Y(n616) );
  OAI22X1 U1813 ( .A0(n570), .A1(n121), .B0(n89), .B1(n122), .Y(n694) );
  OAI22X1 U1814 ( .A0(n557), .A1(n116), .B0(n89), .B1(n117), .Y(n681) );
  OAI22X1 U1815 ( .A0(n542), .A1(n111), .B0(n89), .B1(n112), .Y(n666) );
  OAI22X1 U1816 ( .A0(n529), .A1(n107), .B0(n89), .B1(n108), .Y(n653) );
  OAI22X1 U1817 ( .A0(n516), .A1(n1504), .B0(n89), .B1(n949), .Y(n640) );
  OAI22X1 U1818 ( .A0(n505), .A1(n98), .B0(n89), .B1(n99), .Y(n629) );
  OAI22X1 U1819 ( .A0(n583), .A1(n124), .B0(n89), .B1(n125), .Y(n707) );
  OAI22X1 U1820 ( .A0(n582), .A1(n124), .B0(n88), .B1(n125), .Y(n706) );
  OAI22X1 U1821 ( .A0(n491), .A1(n79), .B0(n88), .B1(n81), .Y(n615) );
  OAI22X1 U1822 ( .A0(n504), .A1(n98), .B0(n88), .B1(n99), .Y(n628) );
  OAI22X1 U1823 ( .A0(n523), .A1(n1504), .B0(n88), .B1(n949), .Y(n647) );
  OAI22X1 U1824 ( .A0(n536), .A1(n107), .B0(n88), .B1(n108), .Y(n660) );
  OAI22X1 U1825 ( .A0(n549), .A1(n111), .B0(n88), .B1(n112), .Y(n673) );
  NAND2X1 U1826 ( .A(n1431), .B(n1433), .Y(n1417) );
  NAND2X2 U1827 ( .A(n1378), .B(n1377), .Y(n1473) );
  NAND4XL U1828 ( .A(n604), .B(n764), .C(n601), .D(n600), .Y(n288) );
  AOI2BB2XL U1829 ( .B0(n601), .B1(n1162), .A0N(n857), .A1N(n1341), .Y(n720)
         );
  OAI22XL U1830 ( .A0(n503), .A1(n98), .B0(n87), .B1(n99), .Y(n627) );
  OAI22X1 U1831 ( .A0(n568), .A1(n858), .B0(n87), .B1(n122), .Y(n692) );
  OAI22X1 U1832 ( .A0(n543), .A1(n859), .B0(n87), .B1(n112), .Y(n667) );
  NAND2XL U1833 ( .A(n601), .B(n1408), .Y(n1387) );
  NAND3X1 U1834 ( .A(n813), .B(n823), .C(n601), .Y(n175) );
  NAND2XL U1835 ( .A(n598), .B(n874), .Y(n1317) );
  NOR2X2 U1836 ( .A(n1330), .B(n1336), .Y(n1082) );
  NAND4XL U1837 ( .A(n763), .B(n765), .C(n602), .D(n603), .Y(n289) );
  OAI22XL U1838 ( .A0(n502), .A1(n98), .B0(n86), .B1(n99), .Y(n626) );
  OAI22X1 U1839 ( .A0(n567), .A1(n121), .B0(n86), .B1(n122), .Y(n691) );
  OAI22X1 U1840 ( .A0(n544), .A1(n111), .B0(n86), .B1(n112), .Y(n668) );
  AOI21XL U1841 ( .A0(N673), .A1(n868), .B0(n763), .Y(n141) );
  NAND2X1 U1842 ( .A(n967), .B(n132), .Y(n84) );
  NAND2X2 U1843 ( .A(n1082), .B(n1081), .Y(n1098) );
  AOI2BB2X1 U1844 ( .B0(n763), .B1(n970), .A0N(n857), .A1N(n1336), .Y(n722) );
  MXI2XL U1845 ( .A(n900), .B(n1305), .S0(n856), .Y(n1307) );
  NOR2X1 U1846 ( .A(n1332), .B(n1392), .Y(n1333) );
  AOI22XL U1847 ( .A0(n182), .A1(err_count[8]), .B0(N813), .B1(n902), .Y(n185)
         );
  XNOR2XL U1848 ( .A(\add_587/carry[8] ), .B(err_count[8]), .Y(N813) );
  OR2XL U1849 ( .A(err_count[8]), .B(\add_587/carry[8] ), .Y(
        \add_587/carry[9] ) );
  INVX1 U1850 ( .A(n1473), .Y(n1428) );
  NOR2XL U1851 ( .A(n1152), .B(sigma16[11]), .Y(n1153) );
  NAND2XL U1852 ( .A(n812), .B(n1386), .Y(n1421) );
  NOR3XL U1853 ( .A(sigma16[11]), .B(n1151), .C(n1152), .Y(n1108) );
  NAND2X2 U1854 ( .A(n1402), .B(n1401), .Y(n1413) );
  NOR2XL U1855 ( .A(n1370), .B(n1313), .Y(n1146) );
  AOI22XL U1856 ( .A0(n182), .A1(err_count[10]), .B0(N815), .B1(n902), .Y(n183) );
  XNOR2XL U1857 ( .A(\add_587/carry[10] ), .B(err_count[10]), .Y(N815) );
  OR2XL U1858 ( .A(err_count[10]), .B(\add_587/carry[10] ), .Y(
        \add_587/carry[11] ) );
  OAI22X1 U1859 ( .A0(n100), .A1(n84), .B0(n500), .B1(n860), .Y(n624) );
  OAI22X1 U1860 ( .A0(n109), .A1(n84), .B0(n533), .B1(n866), .Y(n657) );
  OAI22XL U1861 ( .A0(n113), .A1(n84), .B0(n546), .B1(n111), .Y(n670) );
  OAI22XL U1862 ( .A0(n118), .A1(n84), .B0(n552), .B1(n116), .Y(n676) );
  OAI22XL U1863 ( .A0(n123), .A1(n84), .B0(n565), .B1(n121), .Y(n689) );
  OAI22XL U1864 ( .A0(n129), .A1(n84), .B0(n578), .B1(n124), .Y(n702) );
  OAI22XL U1865 ( .A0(n82), .A1(n84), .B0(n487), .B1(n79), .Y(n611) );
  NAND4XL U1866 ( .A(n133), .B(n134), .C(n135), .D(n136), .Y(n132) );
  NAND2XL U1867 ( .A(n225), .B(n596), .Y(n134) );
  NAND2X4 U1868 ( .A(n1099), .B(n948), .Y(n1103) );
  AOI2BB2X1 U1869 ( .B0(n603), .B1(n1159), .A0N(n857), .A1N(n1330), .Y(n717)
         );
  NAND4X2 U1870 ( .A(n1072), .B(n1071), .C(n1070), .D(n1069), .Y(n1330) );
  AOI22XL U1871 ( .A0(n182), .A1(err_count[7]), .B0(N812), .B1(n902), .Y(n186)
         );
  XNOR2XL U1872 ( .A(\add_587/carry[7] ), .B(err_count[7]), .Y(N812) );
  OR2XL U1873 ( .A(err_count[7]), .B(\add_587/carry[7] ), .Y(
        \add_587/carry[8] ) );
  NAND2X2 U1874 ( .A(n1443), .B(n1454), .Y(n1494) );
  NAND2X1 U1875 ( .A(n1407), .B(n1387), .Y(n1390) );
  OAI2BB1X1 U1876 ( .A0N(n1408), .A1N(n601), .B0(n1407), .Y(n1409) );
  NAND4XL U1877 ( .A(n1330), .B(n1311), .C(n1336), .D(n1327), .Y(n1128) );
  NOR2XL U1878 ( .A(n1434), .B(n1435), .Y(n1438) );
  NOR2XL U1879 ( .A(n871), .B(n1336), .Y(n1337) );
  NAND4X2 U1880 ( .A(n1076), .B(n1075), .C(n1074), .D(n1073), .Y(n1336) );
  OAI22X1 U1881 ( .A0(n113), .A1(n92), .B0(n539), .B1(n859), .Y(n663) );
  OAI22X1 U1882 ( .A0(n123), .A1(n92), .B0(n573), .B1(n858), .Y(n697) );
  OAI22XL U1883 ( .A0(n118), .A1(n92), .B0(n560), .B1(n116), .Y(n684) );
  OAI22XL U1884 ( .A0(n109), .A1(n92), .B0(n526), .B1(n107), .Y(n650) );
  OAI22XL U1885 ( .A0(n129), .A1(n92), .B0(n586), .B1(n124), .Y(n710) );
  OAI22XL U1886 ( .A0(n82), .A1(n92), .B0(n495), .B1(n79), .Y(n619) );
  OAI22XL U1887 ( .A0(n100), .A1(n92), .B0(n508), .B1(n98), .Y(n632) );
  NAND3X1 U1888 ( .A(n595), .B(n814), .C(n225), .Y(n133) );
  NAND3XL U1889 ( .A(n208), .B(n1506), .C(n599), .Y(n135) );
  AOI22XL U1890 ( .A0(n182), .A1(err_count[11]), .B0(N816), .B1(n902), .Y(n181) );
  NAND2XL U1891 ( .A(n1490), .B(n1489), .Y(n1492) );
  XNOR2XL U1892 ( .A(\add_587/carry[11] ), .B(err_count[11]), .Y(N816) );
  OR2XL U1893 ( .A(err_count[11]), .B(\add_587/carry[11] ), .Y(
        \add_587/carry[12] ) );
  NAND2X1 U1894 ( .A(n1396), .B(n1383), .Y(n1386) );
  NAND2X1 U1895 ( .A(n1396), .B(n1383), .Y(n1348) );
  OAI2BB1XL U1896 ( .A0N(n1397), .A1N(n603), .B0(n1396), .Y(n1398) );
  NOR2XL U1897 ( .A(n1393), .B(n871), .Y(n1395) );
  NOR2XL U1898 ( .A(n1330), .B(n1392), .Y(n1331) );
  AOI22XL U1899 ( .A0(n182), .A1(err_count[9]), .B0(N814), .B1(n902), .Y(n184)
         );
  AOI21X1 U1900 ( .A0(n1497), .A1(n1496), .B0(n1495), .Y(n1498) );
  NAND2X1 U1901 ( .A(n1459), .B(n1468), .Y(n1465) );
  XNOR2XL U1902 ( .A(\add_587/carry[9] ), .B(err_count[9]), .Y(N814) );
  NAND2X1 U1903 ( .A(n1473), .B(n1468), .Y(n1496) );
  OR2XL U1904 ( .A(err_count[9]), .B(\add_587/carry[9] ), .Y(
        \add_587/carry[10] ) );
  NAND4XL U1905 ( .A(n839), .B(n1362), .C(n1314), .D(n941), .Y(n1149) );
  OAI21XL U1906 ( .A0(n1444), .A1(n970), .B0(n1445), .Y(n1447) );
  NAND3XL U1907 ( .A(n1445), .B(n811), .C(n1482), .Y(n1448) );
  NAND2XL U1908 ( .A(sig_all_zero), .B(n1340), .Y(n1309) );
  XNOR3X2 U1909 ( .A(n1419), .B(n1452), .C(n1418), .Y(n1420) );
  XOR3X2 U1910 ( .A(n1453), .B(n1471), .C(n1452), .Y(n1468) );
  MXI2XL U1911 ( .A(n596), .B(n1145), .S0(n863), .Y(n1360) );
  MXI2X1 U1912 ( .A(n593), .B(n1108), .S0(n1345), .Y(n1366) );
  NAND2XL U1913 ( .A(n1507), .B(n1331), .Y(n1396) );
  NAND2XL U1914 ( .A(n1337), .B(sig_all_zero), .Y(n1406) );
  INVX8 U1915 ( .A(n1346), .Y(n1345) );
  NAND2X4 U1916 ( .A(n1329), .B(n1328), .Y(n1507) );
  NAND2X4 U1917 ( .A(n1507), .B(n1340), .Y(n1346) );
  NAND2X4 U1918 ( .A(n1424), .B(n1425), .Y(n1452) );
  XNOR2X1 U1919 ( .A(err_count[12]), .B(\add_587/carry[12] ), .Y(N817) );
  OR2X1 U1920 ( .A(err_count[6]), .B(\add_587/carry[6] ), .Y(
        \add_587/carry[7] ) );
  XNOR2X1 U1921 ( .A(\add_587/carry[6] ), .B(err_count[6]), .Y(N811) );
  XNOR2X1 U1922 ( .A(\add_587/carry[5] ), .B(err_count[5]), .Y(N810) );
  OR2X1 U1923 ( .A(count[7]), .B(count[8]), .Y(n1632) );
  AOI21X1 U1924 ( .A0(count[3]), .A1(n952), .B0(n1632), .Y(n1631) );
  AOI31X1 U1925 ( .A0(count[2]), .A1(count[1]), .A2(n952), .B0(count[5]), .Y(
        n1630) );
  OAI2BB2X1 U1926 ( .B0(count[6]), .B1(n1632), .A0N(n1631), .A1N(n1630), .Y(
        n1633) );
  OR3XL U1927 ( .A(count[9]), .B(count[8]), .C(count[7]), .Y(n1634) );
  OR4X1 U1928 ( .A(count[6]), .B(count[5]), .C(n952), .D(n1634), .Y(N266) );
  NAND3X1 U1929 ( .A(count[2]), .B(count[1]), .C(count[3]), .Y(n1636) );
  OR4X1 U1930 ( .A(count[7]), .B(count[6]), .C(count[9]), .D(count[8]), .Y(
        n1635) );
  NOR4BX1 U1931 ( .AN(n1636), .B(n1635), .C(count[5]), .D(n952), .Y(N264) );
  OR3XL U1932 ( .A(count[9]), .B(count[8]), .C(count[7]), .Y(n1638) );
  OR4X1 U1933 ( .A(count[2]), .B(count[1]), .C(n952), .D(count[3]), .Y(n1637)
         );
  OR4X1 U1934 ( .A(count[6]), .B(count[5]), .C(n1638), .D(n1637), .Y(N263) );
  OAI21XL U1935 ( .A0(count[5]), .A1(n952), .B0(count[6]), .Y(n1642) );
  INVX1 U1936 ( .A(count[7]), .Y(n1641) );
  OAI21XL U1937 ( .A0(count[1]), .A1(count[0]), .B0(count[2]), .Y(n1639) );
  NOR4BX1 U1938 ( .AN(n1639), .B(count[7]), .C(count[5]), .D(count[3]), .Y(
        n1640) );
  AOI21X1 U1939 ( .A0(n1642), .A1(n1641), .B0(n1640), .Y(n1643) );
  OR3XL U1940 ( .A(count[9]), .B(count[8]), .C(n1643), .Y(N327) );
endmodule

