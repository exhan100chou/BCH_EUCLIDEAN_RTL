module multiplier_column3_p16(b,P1,P2,P3,P4,P5,P6,P7,P8,
                                P9,P10,P11,P12,P13,P14,P15,P16);

input [12:0]b;
output [12:0]P1,P2,P3,P4,P5,P6,P7,P8,P9,P10,P11,P12,P13,P14,P15,P16; 

//wire[415:0]P;

wire	[207:0]P;

wire BBM1,BBM2,BBM3,BBM4,BBM5,BBM6,BBM7,BBM8,BBM9,BBM10,
BBM11,BBM12,BBM13,BBM14,BBM15,BBM16,BBM17,BBM18,BBM19,BBM20,
BBM21,BBM22,BBM23,BBM24,BBM25,BBM26,BBM27,BBM28,BBM29,BBM30,
BBM31,BBM32,BBM33,BBM34,BBM35,BBM36,BBM37,BBM38,BBM39,BBM40,
BBM41,BBM42,BBM43,BBM44,BBM45,BBM46,BBM47,BBM48,BBM49,BBM50,
BBM51,BBM52,BBM53,BBM54,BBM55,BBM56,BBM57,BBM58,BBM59,BBM60,
BBM61,BBM62,BBM63,BBM64,BBM65,BBM66,BBM67,BBM68,BBM69,BBM70,
BBM71,BBM72,BBM73,BBM74,BBM75,BBM76,BBM77,BBM78,BBM79,BBM80,
BBM81,BBM82,BBM83,BBM84,BBM85,BBM86,BBM87,BBM88,BBM89,BBM90,
BBM91,BBM92,BBM93,BBM94,BBM95,BBM96,BBM97,BBM98,BBM99,BBM100,
BBM101,BBM102,BBM103,BBM104,BBM105,BBM106,BBM107,BBM108,BBM109,BBM110,
BBM111,BBM112,BBM113,BBM114,BBM115,BBM116,BBM117,BBM118,BBM119,BBM120,
BBM121,BBM122,BBM123,BBM124,BBM125,BBM126,BBM127,BBM128,BBM129,BBM130,
BBM131,BBM132,BBM133,BBM134,BBM135,BBM136,BBM137,BBM138,BBM139,BBM140,
BBM141,BBM142,BBM143,BBM144,BBM145,BBM146,BBM147,BBM148,BBM149,BBM150,
BBM151,BBM152,BBM153,BBM154,BBM155,BBM156,BBM157,BBM158,BBM159,BBM160,
BBM161,BBM162,BBM163,BBM164,BBM165,BBM166,BBM167,BBM168,BBM169,BBM170,
BBM171,BBM172,BBM173,BBM174,BBM175,BBM176,BBM177,BBM178,BBM179,BBM180,
BBM181,BBM182,BBM183,BBM184,BBM185,BBM186,BBM187,BBM188,BBM189,BBM190,
BBM191,BBM192,BBM193,BBM194,BBM195,BBM196,BBM197,BBM198,BBM199,BBM200,
BBM201,BBM202,BBM203,BBM204,BBM205,BBM206,BBM207,BBM208,BBM209,BBM210,
BBM211,BBM212,BBM213,BBM214,BBM215
;

assign BBM1=BBM24^b[1]^b[12];
assign BBM2=BBM23^BBM183;
assign BBM3=BBM23^b[2]^b[5];
assign BBM8=BBM41^BBM152;
assign BBM9=BBM36^BBM178;
assign BBM10=BBM24^b[7];
assign BBM15=BBM69^BBM153;
assign BBM17=BBM53^BBM184;
assign BBM18=BBM53^BBM185;
assign BBM19=BBM49^BBM186;
assign BBM23=BBM40^BBM187;
assign BBM24=BBM44^BBM180;
assign BBM26=BBM101^BBM144^b[0];
assign BBM27=BBM79^BBM154;
assign BBM30=BBM92^BBM155;
assign BBM31=BBM68^BBM188;
assign BBM32=BBM67^BBM188;
assign BBM36=BBM60^BBM180;
assign BBM40=BBM62^b[12];
assign BBM41=BBM56^b[6];
assign BBM42=BBM98^BBM192;
assign BBM43=BBM98^BBM190;
assign BBM44=BBM91^BBM193;
assign BBM45=BBM94^BBM175;
assign BBM49=BBM119^BBM156;
assign BBM51=BBM89^BBM191;
assign BBM53=BBM79^BBM181;
assign BBM56=BBM127^BBM194;
assign BBM57=BBM95^b[10];
assign BBM58=BBM127^BBM195;
assign BBM60=BBM99^b[12];
assign BBM62=BBM128^b[9]^b[10];
assign BBM63=BBM87^b[11];
assign BBM64=BBM118^BBM194;
assign BBM65=BBM129^BBM196;
assign BBM67=BBM129^b[4]^b[12];
assign BBM68=BBM141^BBM171^b[0];
assign BBM69=BBM97^b[9];
assign BBM70=BBM128^BBM197;
assign BBM71=BBM130^BBM195;
assign BBM76=BBM123^b[11];
assign BBM77=BBM144^BBM168;
assign BBM78=BBM124^b[8];
assign BBM79=BBM116^b[5];
assign BBM80=BBM156^b[8]^b[12];
assign BBM83=BBM130^b[4];
assign BBM84=BBM160^BBM192;
assign BBM87=BBM131^b[9];
assign BBM89=BBM149^BBM186;
assign BBM90=BBM147^b[7]^b[10];
assign BBM91=BBM111^b[6];
assign BBM92=BBM103^b[0];
assign BBM93=BBM104^b[1];
assign BBM94=BBM148^BBM192;
assign BBM95=BBM157^BBM197;
assign BBM96=BBM151^BBM200;
assign BBM97=BBM159^BBM196;
assign BBM98=BBM110^b[1];
assign BBM99=BBM131^b[11];
assign BBM100=BBM166^BBM169;
assign BBM101=BBM167^BBM170;
assign BBM102=BBM140^b[9];
assign BBM103=BBM148^b[4];
assign BBM104=BBM170^BBM172;
assign BBM105=BBM143^b[6];
assign BBM106=BBM154^b[1];
assign BBM110=BBM143^b[12];
assign BBM111=BBM158^b[8];
assign BBM112=BBM149^b[7];
assign BBM116=BBM144^b[9];
assign BBM117=BBM150^b[4];
assign BBM118=BBM151^b[5];
assign BBM119=BBM142^b[5];
assign BBM123=BBM155^b[5];
assign BBM124=BBM184^BBM185;
assign BBM125=BBM160^b[4];
assign BBM126=BBM172^BBM191;
assign BBM127=BBM176^BBM187;
assign BBM128=BBM169^BBM201;
assign BBM129=BBM153^b[7];
assign BBM130=BBM176^b[2]^b[8];
assign BBM131=BBM185^b[4]^b[8];
assign BBM140=BBM191^b[12];
assign BBM141=BBM166^b[1];
assign BBM142=BBM167^b[2];
assign BBM143=BBM179^b[10];
assign BBM144=BBM174^b[6];
assign BBM147=BBM188^b[11];
assign BBM148=BBM169^b[5];
assign BBM149=BBM193^b[1];
assign BBM150=BBM175^b[12];
assign BBM151=BBM178^b[11];
assign BBM152=BBM179^b[2];
assign BBM153=BBM172^b[1];
assign BBM154=BBM185^b[12];
assign BBM155=BBM183^b[2];
assign BBM156=BBM200^b[0];
assign BBM157=BBM171^b[1];
assign BBM158=BBM166^b[0];
assign BBM159=BBM168^b[4];
assign BBM161=BBM179^b[6];
assign BBM4=b[0]^b[1]^b[2]^b[3]^b[5]^b[6]^b[8]^b[9]^b[10]^b[11]^b[12];
assign BBM5=b[0]^b[1]^b[3]^b[4]^b[6]^b[7]^b[8]^b[9]^b[10]^b[11]^b[12];
assign BBM6=b[0]^b[1]^b[2]^b[4]^b[5]^b[7]^b[8]^b[9]^b[10]^b[11]^b[12];
assign BBM7=b[0]^b[1]^b[2]^b[3]^b[5]^b[6]^b[8]^b[9]^b[10]^b[11]^b[12];
assign BBM11=b[1]^b[2]^b[3]^b[4]^b[6]^b[7]^b[9]^b[10]^b[11]^b[12];
assign BBM12=b[0]^b[2]^b[3]^b[4]^b[5]^b[7]^b[8]^b[10]^b[11]^b[12];
assign BBM13=b[0]^b[2]^b[3]^b[5]^b[6]^b[7]^b[8]^b[9]^b[10]^b[11];
assign BBM14=b[0]^b[2]^b[3]^b[5]^b[6]^b[7]^b[8]^b[9]^b[10]^b[11];
assign BBM16=b[1]^b[3]^b[4]^b[5]^b[6]^b[8]^b[9]^b[11]^b[12];
assign BBM20=b[0]^b[1]^b[3]^b[4]^b[5]^b[6]^b[7]^b[8]^b[9];
assign BBM21=b[1]^b[2]^b[4]^b[5]^b[6]^b[7]^b[8]^b[9]^b[10];
assign BBM22=b[0]^b[1]^b[2]^b[3]^b[4]^b[5]^b[6]^b[11]^b[12];
assign BBM25=b[1]^b[3]^b[4]^b[5]^b[6]^b[8]^b[9]^b[11]^b[12];
assign BBM28=b[0]^b[4]^b[6]^b[7]^b[8]^b[9]^b[11]^b[12];
assign BBM29=b[2]^b[4]^b[5]^b[6]^b[7]^b[9]^b[10]^b[12];
assign BBM33=b[0]^b[2]^b[3]^b[4]^b[5]^b[6]^b[7]^b[8];
assign BBM34=b[0]^b[1]^b[2]^b[3]^b[4]^b[5]^b[10]^b[11];
assign BBM35=b[1]^b[2]^b[3]^b[4]^b[5]^b[6]^b[7]^b[12];
assign BBM37=b[0]^b[4]^b[6]^b[7]^b[8]^b[9]^b[11]^b[12];
assign BBM38=b[0]^b[2]^b[3]^b[4]^b[5]^b[6]^b[7]^b[8];
assign BBM39=b[0]^b[1]^b[2]^b[3]^b[4]^b[5]^b[10]^b[11];
assign BBM46=b[1]^b[3]^b[7]^b[9]^b[10]^b[11]^b[12];
assign BBM47=b[1]^b[5]^b[7]^b[8]^b[9]^b[10]^b[12];
assign BBM48=b[0]^b[2]^b[6]^b[8]^b[9]^b[10]^b[11];
assign BBM50=b[3]^b[5]^b[6]^b[7]^b[8]^b[10]^b[11];
assign BBM52=b[0]^b[1]^b[2]^b[3]^b[4]^b[9]^b[10];
assign BBM54=b[1]^b[3]^b[7]^b[9]^b[10]^b[11]^b[12];
assign BBM55=b[0]^b[2]^b[6]^b[8]^b[9]^b[10]^b[11];
assign BBM59=b[1]^b[2]^b[4]^b[5]^b[10]^b[12];
assign BBM61=b[0]^b[1]^b[3]^b[4]^b[9]^b[11];
assign BBM66=b[2]^b[4]^b[8]^b[10]^b[11]^b[12];
assign BBM72=b[0]^b[1]^b[2]^b[7]^b[8]^b[12];
assign BBM73=b[0]^b[1]^b[2]^b[3]^b[8]^b[9];
assign BBM74=b[1]^b[2]^b[4]^b[5]^b[10]^b[12];
assign BBM75=b[2]^b[4]^b[8]^b[10]^b[11]^b[12];
assign BBM81=b[2]^b[3]^b[5]^b[6]^b[11];
assign BBM82=b[3]^b[4]^b[6]^b[7]^b[12];
assign BBM85=b[0]^b[2]^b[3]^b[8]^b[10];
assign BBM86=b[0]^b[1]^b[6]^b[8]^b[12];
assign BBM88=b[3]^b[5]^b[9]^b[11]^b[12];
assign BBM107=b[7]^b[8]^b[10]^b[11];
assign BBM108=b[8]^b[9]^b[11]^b[12];
assign BBM109=b[0]^b[9]^b[10]^b[12];
assign BBM113=b[4]^b[5]^b[7]^b[8];
assign BBM114=b[5]^b[6]^b[8]^b[9];
assign BBM115=b[6]^b[7]^b[9]^b[10];
assign BBM120=b[1]^b[2]^b[7]^b[9];
assign BBM121=b[4]^b[6]^b[10]^b[12];
assign BBM122=b[0]^b[5]^b[7]^b[11];
assign BBM132=b[4]^b[5]^b[7]^b[8];
assign BBM133=b[7]^b[8]^b[10]^b[11];
assign BBM134=b[8]^b[9]^b[11]^b[12];
assign BBM135=b[5]^b[6]^b[8]^b[9];
assign BBM136=b[1]^b[2]^b[7]^b[9];
assign BBM137=b[4]^b[5]^b[7]^b[8];
assign BBM138=b[4]^b[6]^b[10]^b[12];
assign BBM139=b[0]^b[5]^b[7]^b[11];
assign BBM145=b[1]^b[10]^b[11];
assign BBM146=b[2]^b[11]^b[12];
assign BBM160=b[5]^b[9]^b[12];
assign BBM162=b[5]^b[7]^b[8];
assign BBM163=b[0]^b[7]^b[11];
assign BBM164=b[1]^b[10]^b[11];
assign BBM165=b[2]^b[11]^b[12];
assign BBM166=b[10]^b[11];
assign BBM167=b[11]^b[12];
assign BBM168=b[3]^b[12];
assign BBM169=b[7]^b[8];
assign BBM170=b[8]^b[9];
assign BBM171=b[4]^b[5];
assign BBM172=b[5]^b[6];
assign BBM173=b[3]^b[12];
assign BBM174=b[4]^b[7];
assign BBM175=b[6]^b[10];
assign BBM176=b[1]^b[3];
assign BBM177=b[4]^b[6];
assign BBM178=b[0]^b[7];
assign BBM179=b[7]^b[9];
assign BBM180=b[3]^b[5];
assign BBM181=b[1]^b[8];
assign BBM182=b[6]^b[9];
assign BBM183=b[3]^b[6];
assign BBM184=b[0]^b[3];
assign BBM185=b[2]^b[10];
assign BBM186=b[3]^b[4];
assign BBM187=b[4]^b[11];
assign BBM188=b[2]^b[3];
assign BBM189=b[3]^b[5];
assign BBM190=b[5]^b[8];
assign BBM191=b[0]^b[10];
assign BBM192=b[3]^b[11];
assign BBM193=b[2]^b[9];
assign BBM194=b[10]^b[12];
assign BBM195=b[0]^b[9];
assign BBM196=b[8]^b[11];
assign BBM197=b[2]^b[12];
assign BBM198=b[6]^b[7];
assign BBM199=b[3]^b[11];
assign BBM200=b[1]^b[6];
assign BBM201=b[0]^b[1];
assign BBM202=b[2]^b[3];
assign BBM203=b[2]^b[10];
assign BBM204=b[7]^b[8];
assign BBM205=b[10]^b[12];
assign BBM206=b[7]^b[9];
assign BBM207=b[0]^b[11];
assign BBM208=b[10]^b[11];
assign BBM209=b[11]^b[12];
assign BBM210=b[3]^b[12];
assign BBM211=b[7]^b[8];
assign BBM212=b[2]^b[10];
assign BBM213=b[3]^b[11];
assign BBM214=b[10]^b[12];
assign BBM215=b[10];
assign P[1]=BBM166;
assign P[2]=BBM167;
assign P[3]=BBM140;
assign P[4]=BBM141;
assign P[5]=BBM142;
assign P[6]=BBM168;
assign P[14]=BBM169;
assign P[15]=BBM170;
assign P[16]=BBM143;
assign P[17]=BBM100;
assign P[18]=BBM101;
assign P[19]=BBM102;
assign P[20]=BBM141;
assign P[21]=BBM142;
assign P[22]=BBM168;
assign P[27]=BBM171;
assign P[28]=BBM172;
assign P[29]=BBM144;
assign P[30]=BBM103;
assign P[31]=BBM104;
assign P[32]=BBM105;
assign P[33]=BBM100;
assign P[34]=BBM101;
assign P[35]=BBM102;
assign P[36]=BBM141;
assign P[37]=BBM142;
assign P[38]=BBM168;
assign P[39]=BBM141;
assign P[40]=BBM106;
assign P[41]=BBM147;
assign P[42]=BBM56;
assign P[43]=BBM57;
assign P[44]=BBM76;
assign P[45]=BBM77;
assign P[46]=BBM103;
assign P[47]=BBM104;
assign P[48]=BBM105;
assign P[49]=BBM100;
assign P[50]=BBM101;
assign P[51]=BBM102;
assign P[52]=BBM100;
assign P[53]=BBM110;
assign P[54]=BBM111;
assign P[55]=BBM40;
assign P[56]=BBM112;
assign P[57]=BBM78;
assign P[58]=BBM58;
assign P[59]=BBM57;
assign P[60]=BBM76;
assign P[61]=BBM77;
assign P[62]=BBM103;
assign P[63]=BBM104;
assign P[64]=BBM105;
assign P[65]=BBM103;
assign P[66]=BBM116;
assign P[67]=BBM148^b[10];
assign P[68]=BBM79^b[11];
assign P[69]=BBM117;
assign P[70]=BBM118;
assign P[71]=BBM80;
assign P[72]=BBM112;
assign P[73]=BBM78;
assign P[74]=BBM58;
assign P[75]=BBM57;
assign P[76]=BBM76;
assign P[77]=BBM77;
assign P[78]=BBM57;
assign P[79]=BBM41;
assign P[80]=BBM119^BBM174;
assign P[81]=BBM83^BBM175;
assign P[82]=BBM42;
assign P[83]=BBM60;
assign P[84]=BBM84;
assign P[85]=BBM117;
assign P[86]=BBM118;
assign P[87]=BBM80;
assign P[88]=BBM112;
assign P[89]=BBM78;
assign P[90]=BBM58;
assign P[91]=BBM112;
assign P[92]=BBM62^b[3];
assign P[93]=BBM63^b[1];
assign P[94]=BBM64^BBM176;
assign P[95]=BBM26;
assign P[96]=BBM43;
assign P[97]=BBM44;
assign P[98]=BBM42;
assign P[99]=BBM60;
assign P[100]=BBM84;
assign P[101]=BBM117;
assign P[102]=BBM118;
assign P[103]=BBM80;
assign P[104]=BBM117;
assign P[105]=BBM64^BBM177;
assign P[106]=BBM65^b[12];
assign P[107]=BBM87^BBM178;
assign P[108]=BBM15;
assign P[109]=BBM27;
assign P[110]=BBM45;
assign P[111]=BBM26;
assign P[112]=BBM43;
assign P[113]=BBM44;
assign P[114]=BBM42;
assign P[115]=BBM60;
assign P[116]=BBM84;
assign P[117]=BBM42;
assign P[118]=BBM83^BBM179;
assign P[119]=BBM87^BBM180;
assign P[120]=BBM67;
assign P[121]=BBM1;
assign P[122]=BBM8;
assign P[123]=BBM9;
assign P[124]=BBM15;
assign P[125]=BBM27;
assign P[126]=BBM45;
assign P[127]=BBM26;
assign P[128]=BBM43;
assign P[129]=BBM44;
assign P[130]=BBM26;
assign P[131]=BBM68^b[6];
assign P[132]=BBM49^b[7];
assign P[133]=BBM89^b[11];
assign P[134]=BBM10;
assign P[135]=BBM2;
assign P[136]=BBM3;
assign P[137]=BBM1;
assign P[138]=BBM8;
assign P[139]=BBM9;
assign P[140]=BBM15;
assign P[141]=BBM27;
assign P[142]=BBM45;
assign P[143]=BBM15;
assign P[144]=BBM90^BBM181;
assign P[145]=BBM69^b[2];
assign P[146]=BBM91^b[1];
assign P[147]=BBM30;
assign P[148]=BBM17;
assign P[149]=BBM18;
assign P[150]=BBM10;
assign P[151]=BBM2;
assign P[152]=BBM3;
assign P[153]=BBM1;
assign P[154]=BBM8;
assign P[155]=BBM9;
assign P[156]=BBM1;
assign P[157]=BBM92;
assign P[158]=BBM93^b[0];
assign P[159]=BBM94^b[12];
assign P[160]=BBM31;
assign P[161]=BBM19;
assign P[162]=BBM32;
assign P[163]=BBM30;
assign P[164]=BBM17;
assign P[165]=BBM18;
assign P[166]=BBM10;
assign P[167]=BBM2;
assign P[168]=BBM3;
assign P[169]=BBM10;
assign P[170]=BBM95;
assign P[171]=BBM123;
assign P[172]=BBM63^b[0]^b[5];
assign P[173]=BBM70;
assign P[174]=BBM71;
assign P[175]=BBM51;
assign P[176]=BBM31;
assign P[177]=BBM19;
assign P[178]=BBM32;
assign P[179]=BBM30;
assign P[180]=BBM17;
assign P[181]=BBM18;
assign P[182]=BBM30;
assign P[183]=BBM149;
assign P[184]=BBM124;
assign P[185]=BBM65^b[2];
assign P[186]=BBM125;
assign P[187]=BBM126;
assign P[188]=BBM96;
assign P[189]=BBM70;
assign P[190]=BBM71;
assign P[191]=BBM51;
assign P[192]=BBM31;
assign P[193]=BBM19;
assign P[194]=BBM32;
assign P[195]=BBM31;
assign P[196]=BBM150;
assign P[197]=BBM151;
assign P[198]=BBM36;
assign P[199]=BBM106^BBM182;
assign P[200]=BBM90;
assign P[201]=BBM97;
assign P[202]=BBM125;
assign P[203]=BBM126;
assign P[204]=BBM96;
assign P[205]=BBM70;
assign P[206]=BBM71;
assign P[207]=BBM51;
assign P[0]=b[10];
assign P[7]=b[4];
assign P[8]=b[5];
assign P[9]=b[6];
assign P[10]=b[7];
assign P[11]=b[8];
assign P[12]=b[9];
assign P[13]=b[7];
assign P[23]=b[4];
assign P[24]=b[5];
assign P[25]=b[6];
assign P[26]=b[4];



assign P1[12:0]=P[12:0];
assign P2[12:0]=P[25:13];
assign P3[12:0]=P[38:26];
assign P4[12:0]=P[51:39];
assign P5[12:0]=P[64:52];
assign P6[12:0]=P[77:65];
assign P7[12:0]=P[90:78];
assign P8[12:0]=P[103:91];
assign P9[12:0]=P[116:104];
assign P10[12:0]=P[129:117];
assign P11[12:0]=P[142:130];
assign P12[12:0]=P[155:143];
assign P13[12:0]=P[168:156];
assign P14[12:0]=P[181:169];
assign P15[12:0]=P[194:182];
assign P16[12:0]=P[207:195];










endmodule
